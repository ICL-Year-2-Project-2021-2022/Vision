��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	q�v�Z��\R�w�0xtʎ5x5�������v�7\M�k���%n;c-<�<;�`.���B1�7���[�D�\�A��fIj�)����懋�f�7`_�%�E�i�j��yF���^�s�[wg`}vёp�M�=&d.�ȩ$7l	�$����>&R=�M� N=;5k�B���t��7�@>j�c�� �������P�����8��Լ����Y-%(Q�"�{�-�y��< }
��_�E`F���o��)��i�+o��]�KD�(<�~
f�(�Mo�^A(�����8�Bٱ�4Ou�:������/�M�f�(�����//�|�.��&�l*]��?�v��:>k�r�� P���'���#^yĥ���\�t��p�>cY}��Ƃ�	�	�B�٥��V6$�1q���<=�L,���TA�$�{Q�����Ee���νẑ*aD���!ռ	�s���e`�'�00��:^���(t3QV�"�|Q�w��X��\:i!�6�����M�;6���5��Y��uJ����Rey��F��M��d�ua�A7��K��[�4�'F8��0�ѣ���q
��@�ʸ_⿧=,�0��p�����VB�w~  mq�͈V�*���Q��P�iJ�)��\+�S���ԏ�gʥ�U2�����!�Z5i�7/�pGO��\ԅ��4<�ٟ�phCd����0�eP=W�EA)�T���_ ��gs�	A�oz���<Q��0V��b�"��qee�� �w�o|�<������2.�>>� J�����&�ڒ�a�<G�S]5C3�,vj��m&��H�����)��0"n��S�
�(��Т�>��g�����/����4l��������Ra0Q=Q�x�l�@�rt
�Z٪���׆�f��Z���Z��G�>��	bY��f�MZ[@t!R:a�u|3�6�����s����owaKx����ĳ�舻��XA[:�;��:ѯ��5�i��y��ⴂ3|轪l�k�%,���}��`tXl ������F�r�����K��g@�!)���v�2.張����3C���!NxZ�\/�7�:��Zs��dkl�lܫĴ�V���u���獵��ʠ��s�� ���O���H�������u�&ƆV��%z�&�}�=�	ߕ���$��~ӛ0��XX߫�P�����ĉG�����;u�7:&���`���Â�|�E�����[�����x���Յ��{I�Mg��B��ဥo ۸$觊�21X��&%��g��ȖfE-/57��Y�h�A�4[����x�֝h��|�o\��$���	ć9W�%<b7QUr���8�妧��V+��O�=�z�s �vA頱����ht܉���{P�L�;�ć�?{�$�Afk>{��^���@�\:Hj@�~��4	u�u8KÌ-���-vg��L�)Zv�26����O׎04H�Kbj�j5dyA.Z�-ac&¸�Q��E��ژ1>=�7KgG�]�j#Z��el���O7�'gZ���\����_�s���P���y��ǨrV*���3�M8R,%=]�����-�yAT�Z�	ݝԑP���	����t(���9G��5���M��	=�7�u�,�B�k����QT0c{I۽���8�F
�,���z=����󷄗i�����v!d
s�{�_ ��rT�_Fڳ{����G�eu���r�C
7Ϊ��f&�cX�i������&����1��b���W��s�&yYL�n��.�h����1kG�'C�45���B��{Uwt�+����ެ~�v�O㗾��I��R��R E��mD������9G*�la��u�;r��Lyi.�oX�Vt'T�8�yKW�"���E�:l������n��`K���Z�݁���0�w���-!��\]g��'�� &k��@�g	HF���ѠK����X�C"U�Y�m@ޔ�ჩNҏ��1N�ؗ}���5�%�'B��:b)��^Em9�c�}f�3��3����c��^�CBe �g��X!�,1�l�a~$�{�rB��W�K�s����y��z�ȢM$�՞L���%1b<��i��L�u��	�I�Y��qv�,�>UՅ��A>`�n:��7F>��&�-e.�s�`�M���^O�@c�� �L���h/{�g�^���3��_aˌfJ6�!��Bȷ����k��H�F����)��� YR
Y\`�Q��W8St(�|\Dm���=R�#FO2i^�G�����kU)TåƯ���i,�@��|��ٱ[T@��M���c�A�9C�e=���r{2��v4i���1�Ҋ�=�V�f��;�	�O&��͛�Nmꚽ���(Wy���6=�I:X&�{'\�������\ג�E.�&�g'S���s-�m:?�A{k��"�/K�P]�s��@6���������"�\5�K���3��tT��+�}�j�Jw����,H��d� �6��[�}��� ���0bT�l$h';l�݄���zo�bJH�'�-�t��ɋ��N�ŗ}.I��t�C����"�qcq��'*�h,Юㄦq4��m�����c�S�P)
�\��~�6村�>^�j&�\�+&G�=��	�wfx?j����icIι��	}�c��D�7��ľ��6eg>\ �u^7y�H��%-/�Ut�MF����\M-Թw��r�����q�,w�=��5�IA���no�� G� %����J'�+�T(j�҅��)[HnY�T��B84�9��ke��t����f��[%j��p�2�:��	#�t\P�Ňp��&p�Րf뫡7!i��ık�7@o�X�ݛ�f��︓ShB�͒���㔀�s��� *kN��%X4V�K� �'o���$��B�ŝ+�DG���	��)�2����l8Ppl
S�'8n��
���9�ݩ`���XC�vn�ph��G�pl�ϙW��e�Nll흯SZr<�[�P���B�ZD�Je���ȗ>A��7~��D�̒]s��5,U���Ζ��c~������w�}��Jwt�`g%��)��������ɍ-��f��UQxE��S�?+�ų>��8�\a�=�LQ�H��!��{r�fE��=Uw�Q�דϽ������9U�R���B��LL����#C�Dp�/9��t�Q0��FG���!W�on��a�A�30% ��������%�V8��(�p��aO2[�����` ���´�O%���k�ؕ��,�~~�xˑI��H��՘o-,����eƚ�ڣv��̾�v,�	��Ԅ�Mٚ��t�����%錂u����C��K�8��[T�S6@-8?��\1=��`�x&/I3��Mɤx�L�ϑ�	^.z���n��LXy��V�)��I2j��H9x�:�h�A�	)�o��4Ƣ�F5����2���j��a����A-�1�"&�n�OK;,�&X4bn�=JB�D���b/,_��wv�G�ќȉ��"�&���!��Ў����h���Gq!�����FP?m-��2��8H��z����u���B{�)$��9ZJ���u���k���$�Y��L����� a�#�N.��-�t�{�W��.Y%�����j6��ݡHx��NI9�<��y+ɶE��Ɣ$x���a"z���4�~M7N)�t{3�ۺ|�B��_5F�Ylis#��ܖ��~�T�Qr]��Fb/�J|d�g���'`u�r �|��}��d�ժr!�F6!AJ"�|�q��ᚔF�U�)�|A��&��[��y�v��p���ׁ�JD쓝VIwz�z�$ �^`I5h#u�a��T͌*g&�&^{��ͽ�?�h�}���@�Á2�@R��'s��_�zS���K��$.�T�y�}F
�d?��" �~�BA@��ۻʡ���̚r>���F�l�!��gv$x��:�ۼƙ��_x�q�U�%(�8j���}ODC��D҆����)a���5�p߉�M��x�yIt9��KJ�e<��m��;����2�%��;����	Eʭ�(�k�w�9(���Q����Z� F�ЭR�=��0.��!)��0��xd%�:�U�Z�����4�1�Ji�W'�3�.��*�e�oB���߬Y	�m�՗3EV�>��n�a�ɤB��=��Hɭ�*�}.�-`Æ#��ܿl�K}	v8b�e��m$��d��tH���$�njm����LNV�n@ bQ�/9^�����k�p�y��d��K��ط�5����-	ѧ2'�g���sq@���s�,�v�V�l�xX�~�{G#��ȩk}3�<2�KS߆��$��`�����Đ��?0F��M��Z���ھ�N/9:/t�
.��.�ѡ$�B4�;[����k�1���(�p%�R�T�G+&�;w*wW�j{PU��-��9�<��E52:��t�F>[�g��0�P�E�`��T!1�������gV�yxO���#;d��JhN�4�o�����n*�=�ďvN����E�7B�9��A�ӵ[�!��L�P\��/Ŵ�����xcq�D���P7��R�&�a����24��	3�/3��5��`�L{I����!B���c�^�[o����KI�]�� �K����,�� !�G��?�8�/�{.���yD�PebB~JU{	X�#�ڒ�y�IoP�&�ӳ����mm&U3JK�L��@�~��@�h��C���gd%r�^'Ӫ2��q�c��#9�L�-$4z	˩���>F�+�R��l]�I�Q7z���(�+'�a{B�^%zpA8�Ґ�0R�k��I��[J���21{�|�3��}F�8lk��=՚�3٣����X��f�W��hSNA�����H�!j���1��"���fkx�K�ԩ;��*A��:�J�uL�I�'vh3���*������ O�Gν�B�7/!&I���V>�����z��+^Y��0?)m5(]�9�#�}_�.ݡ3�L|�0�L
R���=��@fYL��6k�&]z!j�38��Q�K��^#ٞݚc���kM43�l��grj|���J�V�f�H���$���p pFÚ��z��f�!>_}Z�V�����"C�E���
�w;�ĺ��f4��� �������Y?�L?��݃��֟��Q�ԓ���né���"�n���is��K^̚~���lZ�Ϋ��g���+�!�⃩�FG��;&���l6��㠡�(�c�"<�V�T�Y���p��lt���ɜ���-�����'U�`9���@m���
Lq����&�d֪�|1+֘	󦥁D?�i3�CYG&�O��_E	�kq��������u_�i�=l���W��{jJ������NLQa'q攽�Ճp��G(��&�;���$��/�9�!���p���rXW=7L����%t<��Lٞ��I�N��O�/7�G��щ|��Ws���{ɏ������V�GLp�n������2p�p��|L�X �;�gV�WQ@���~t�]\>f�����!�,�+׍���ك�NN����"� ��g�{�bC�4���B>V��Hgym��7<��P`%�M.\�8�=?)5��'k=�v�(�������B��Y
X����Z?��(1I����lp^9A�/����,?�nI6�������N7!��� ���Ǘ���-(0<����m����P�5m��L�L&��8���B��gKim$���]��-��L�[�L�F�H�z��8����,��6�K-ĩ�����G��=���L0Ut	�.�:>�ߤ���>���G�`�P/�.�EWij��8�]�ׇ����b,�R�n�83z�%Ө�S"�#�|�V����@��-���8�xq�`�2��K�K�靿8�8�@�s`�}�*�����A=�p���d�m��e��p��`�O���9%���{2���m��*(xU^QT�f�V�G*�{��I��p���Q3v.ڢ��~/�X~G�4<���zR���Ζ<XQ���޼)�y"[�a[`��f��
;|1�O��k9�pu��ʴ��o�9	Ͼ�rW�k��Տ���
<�����3��� ����������
�Wڢ#�b����cلo�������C�0�h�&J�S�����q	��.E�v`�_L��\�o���i�6Fى�>�Gm*�}�x>�ɟK��q��塍��Ǜ~oѝ��x��,yASjx��� pX9���ND]�&�đ�?P�y�f�G�Y=��L��)�+Of1�xU�����
�44�c�/�ga�_dؖz�+.w��3��=�nŹn�A���f�lj�֕t�0%Y���w���3�`
��*�ܫE'	���]]�8��䛙���.%^f�je��� 9��8>ӂFIhZa=k����ڐ�w}[3�C<f�.&Bc�n^�ʍ�����V=��n�E�qw��66�Fa�K��ry>#}�S���?���y�2`�����{㡨γg�ʙ�KeE�gO2��3Ⱦsގ������v4��:`:�:L�7�.�(��@rpO;�!���?��N7pܯ��*�1��c��Y_Π~�B�)���z�n^��Z�b���}w���R4�t�T����h7f�f�Q�R+���y�T��c>a��0���䤭R�Y��CG�BS��ְ^LG������5��F���'�>@+2j�� i�&����1�	m�+�e��%�3�aЁ�l&��9t�ǚ!��qڌ4�{02U���}m�b����mz�J�Gy��0�� S���ptް:�̽'��U� G�8�YئP��*�l���;9ӅM�C��~
���:W���T�L�l*��d��V����֏D�D��lʪs����C�[�<���b|��h�����"�v�g��jL#)ن� +s�i�S����t����ג���Cm��N�nv��
�zj��X�Kq�♜`�$7�Sߕi@h�Y��}������c�ۆo�H-�-6*��F�wA�w����FB��륦�3&5��b�+]x��Q�i�����W�9�pe(#���Di�%R�P���I�#�T�}�>�3xqk�h>�����B�$K:�e�.�.�{OCD9�2/S�R��Wg�7{ȵ|��������>K�a����\5�r޺@J�Gw�K���t*'�Q.P�尪5
V�?���A��?D��^�9<�cH?L���\�C�r7a��o�m����Q("����.��@]���(�z]������8N���3�3XXք����:鸬a7�Q�����ɘ���g`.���k��ܱMx�	�S)��˔�5.���i�e����/z��2`*M/��>u��8I��^�.|�a)��?r��lC����]�"��;�MsS��s(�B�����,%���C%�S�%1mԭ��x�!-Nt�h�I$�.Z5��Q�X��ya�@��k�> (��3*e���(c����rd����R5o&a�k�{�@����,�f�=ϕ<���MO1����aO�x��:vFk+il6/�ꆄ �_j�i��~L<��k:F��@s�h<r��(�Bc��d;[q"��_2�R_
�o�#�/z��)`�p
ao�VwRu�)�Պ���)#Q��4�}��y��1�t�rf���_r���|/f�3C�C�Aw��")Ӱ�?�U��A>�b��W<�_�*���)���27)���Z�w�0� �ōe�s
벰9"���L�=U�v~��n����n�<�l8]�npx�~���Nr �0���X6UK/f��_�|����4��w�M+r�=�(�^���E=�ay[�|îw&��r6�B莁ei6�e���{��9Q������p�!n �{����7d�� Z��Y�����vʓ{��=bt=#Q���I�=�'
I2b�pQO�#�ы�� ��+`imWb�"p�/'ݡ����g���(�݊��8�j��x?}.�oKl���y^V�}��쬵�����q+�T�1�����n�>���NO�P�<�u�v������=��<���3<7n���36����g�+���zM�7cB���YՓ���3��f��#(`n>�r-�^{�c�=*��k %�O��Z�<�H@�PE��rz��?^������S����K;*!�{f���[r�-1-��kT�w�]��ݼ��q"�u�-	t�e]P�\s ��+�1i1T-��]����U��KLEy�l�rځ�P�ܔ�����
���z-L���B?��,[R�z�dX�N��#y�n�ǃY��0��P�������7ٞ�c�Ae�Ze��Ӕ�n��*i��e\��w�K�i=�Ľߍ�+v�ٹ�����/��gA�h+�焐���"=��ZO�[��1��<N`(�tG	�{S��j�(�n%�XZ)��hiM"KG���(����R��}��vٽ��>1M��ƽ0�T�t��(�`׊y�RX���7ps*Z�9iU
�<�����]m,�PA�PE�ʾ(0����	�|K��tx���$�s/���>Ucl/����g�������'+"��[��/�!Ik�"'ȁ�n�ћT�`hN��;F������޴)��r2-����]�&����f ����ct����C�z�n�Z�x8�S���ٲ4��������E��_�*<N��?bR"q��#K5b�,(�b��D�0G.vd��Ƌuz�K�2wPTϢ�	�~��z�R��=���Ƿ%��<L+��H�dW�E|1Ӝ��K��d�Y������xs�i�۶B.V�m�ѿ6=��W:R/SC����QNj̻\t?���K�Jވ�������fYC� ��X��x^G�n��4 ���B6:��I��2^�A���7VF���`e�54o�i��6��z#����D������^�P��`�Iz�.�5���I_�G�qMgt���ŗخ�wkCGL�
5�,�cP����ҦO�7�GY��:oWhm6�Sxk`@��.��N�"�9 ;�Ɯ���&�`�}��
|8��������XT�'0f�H4�WU����K������4,fn��{�<S���S��|Z$W�.ok�2d��jw��?q�����?'��e�:G���� �W�F���8���X|���O~&�
�|*@����񃆁t�G�@���n8���J��l	�}Ԗn��������VF6�!Z�ƥ$�e��y_S��&��+f#��o���5:8aQ��ܐ��
`�� ڒn&5��b���`1QyE�[�YJ|B���T�˛�4G��s*�ц��0k�����7��p� {3_�q�m���>�w��@�e���p.>q+�����ě���2>��ⷋV5u��Fo!6�Ȑ� ,6���p����'M-��E"�y�9�s�]��@���@r��:���lڴ�zcF"/6At���8n�&|hQ�ر�*sf����I��]Lsv��A��q�2�AO��ɵ��=XzN���j\�F��6�ilR˴J�#m�cv�O�7�N�C���b_i�4�ń�2L2s���8r2�2������)o�Lg�KC����H�p���h���kriᘪ�Z:���hu%��YDP�� 0|�	4lP�z)�����>)�_hԇ��L�7���br5w�6aP�R:ܡR3y/�m�n%��"���ti�*c�Z�vV!��?����<����Cퟌq䅄_�z��<����$����x#��F_��a����NT�*��Y(���#%�ŢÇ����t���z�`�}�t�&�.	��lP</};�����#����S��!ψhq<��'d%�o�'df)��d6W+PEr�*"[����{NlGQ!�[z���Q|���̬7��J+�Y%�\yw�J�e�47 ��r�A�Z��Tl3U��ٙ���X蹪+��P��s05�z\Xó{kK��_�C� w�e���;
�Su!b�J{��,ī�-(� �ՐX��ɼ�Xtf�#��Q�&w�����%Ez��!6J��|�ڂ���}y���r5y�y&������`�i����n�0��[���K��Ԡ�J��%&���(�0��zp�5�t��t�,���d	\�Z_#bN�e>��z�NI�2ؙ�f�=����t�� >ٷ�̖�i�x��ME��ҩ\��0Yq�Ʃ��[�V����􄸢/\�� ����op��S�N�=1��c�����ӯm���B�����S��H~�ZG�ݶPϾE��`O�f�/|�'�ǐ� ���Ejp�N�U�J�%W�Y)�^TI����/g`*��%a�̵�n�*nj��oG��4�:�T1`��	F{0A&�O�$��\dz�~Y;�,��$��3g=8Zoi���Ug��y��cJ�ˮ�'G��'�ui\�{����ӣ3����E��EΪ ���+�����v���vG��ׁ�y� ���u��������FO��.Ƨ;�O5���dw%���A��=�(~��X���[����Z�K�so$H+ u�;q�&ѨHN�����n@���x�	�h4�㍚��5�D���X�P$��;�T`�ai��CK��v�	����� ������/��-�ad���C�wg�Z͍�@"�K�k>��
���L���!b�B��k�d9h���ABę�j��l��G��zBJð����X�ȱ&��F����co��6R� �g�h�_w�����̆���`'$łĽ�݈Ssѥ�b����
��yQr�?�0����!3�k`�e
/�l�^�5�!�ѷ�b}��d���-װ{��|�ڶf�b[N���&��R�#��&el"N[�GH* ���AQ���+0&S���4SW��%c��������?��r� �G��,!;+~��j9ѕQ/)C�2 n�ʪ�v�feA(	�[���a��V=�E�^�4�ϞZ��[�ڠ1���ݻ���Z��t���\��RA ��^���6������b���>�h��L,r�-X�ً�����G<]��������BZ�t�w?ͯG���9��OS�f���t=��	E�%��]�$x��w�K��KB�*�;���]�����`�ҥ��7�(��������D��G_o�L+HI��Ԟ�JϨꯇ�23�K|��s��#ٯ�}3D�6]?�np{��]�c�����v? ��I�r�}��r�D޽Mrur��W���:M�ܽۈ��tICkI��_�����9Y-���~�6C_"s�|���Y��˪?�H'��0�b|�z�G/��"Z��+Ț�s���m�.�U��/s�G���?�;�siT�=+�U9�'6x�������;dFW�N-3.z3A#^�l�9�D�Å�{���UUJ6H�,b9�6GA>��F���]]��=�V,�Czl��� ��ɜ����rBo�T.�<i��0\���$lh�����`��K���3�>����èh#R3�'0U~��$_�_�z|�;~}(	h�{>U� IDD`q�[�ˁ�`�ܶ�g�t�4�w曒��Dc�hceGb8��U`)M�hrTV�j�"p�x�El�xD�1��Y��t��k0oI�ez����;�J]DH58ƃ��w��c�ȍYo5�:sNC��^�U�L�s�#��R�.���L��t�nD�G�;H��F�����C(�zj LkO�@ڂ���������]��#�F8�6�پ��������/��bd�~�='�~�9|zo��z#�4�g���0i�-�ރ� �e�2��(��<lɗ`5��kz�1����#AJ�۽+���%KGMv�/tt���S/坿h�n�K�GH����x �~��>B#�y�p>�1�fu����4 ��B0�4��ȃ�ͣ��~�!�	Á5~�^eE�{�i�.|3�$�%7���m�e�yr�0b����31S������^�
�ek�5~��g�9e�[��f]t�)�U߳z�d�z�ԶV~,�f���Ԣ!�	���[����ܩC���?u�X���-�9���%O:�!�8̚��O����6�vi���Ed��-������#��u�o�.+%���fq�E�ScW|��\�a*��\���/�����pLy_���|�{7x���X6���YB��5����(\r������>r�Z)�V�U��R���DN�]����z8Q����o5eO���.�`&�b�qC��X%�Rl_7����9+V����^T�o�+T�t�7*���蝐��(��=$f'n�m�Z�cAJD��`2U��i[�N5@F��k[o#AD�$tl�QB��ug�rw7���F@�?L�_-��nv1 )/�����d[�-0���^�����k�d=Mdp�#�qs�_��?'r/���n�Y7���.��u�����x�������I =;G�<LD�p�G�7܂��"ע_��%e���Ic�8��ߛ[fb��Xy#ۿ��o4G��d�	���Bn�`:�nB��_�ƹI���@�oX-9�-��Ę�xg[Y�R�=�( �͈��B��\wH}W���"m+� =I��ٷS�`��*��3'9A��S�>�|�옘ȋ��i+���{]ު10�������k����m=��6�
��Á�o��=��,�D�}"�5?|�\�jpQ���z:#�l���"۪��fŨl�^[5�-��N��/z��Q����F��R`iX9�T\�}�G3Qo�WVuڳN�D��`ÏY�@�Nq��c�n��� �,��I�A��6h��@�5��GEE�/�e��1�����>����������+��q�+����݅�O_Ӽ*��0r��Ӄ����Ija6?+d(Hƒ8p�7M�~	�� ��[3�]�����T�O)L��N��T�IW��~���x"�!���@x$�Jmۢ��=5�i�r�J)���*�`A�E������F���9�n7�뉼A̽�5P�i�+��^/*��4n|}C:�&�_vC��O^i�yТӏ�z�2��hc)l1�5�cҿ^������W��g�%�0�$�|8�K��@C�^��p�Jqm��0�ᩂ�.����P=<�I���v�mek!d�e�Kܚ��}�W}����Դ9��o�aG8M�c*cZF�-s<'��W���nH�+�������	�FKAbKփ<�Gf�m�K1����S��FJ���Z�𛪓�/\��1�)���s�6+�/b!��L)�@��%/ZXm�n~$~t�W�&"e����M�A��̇욋����n�Wmk�T~�#�� ��U���)ڨ�D�|s��/��@Т��L�)x_�6dj���U����	G���ϟ8��/�à�N�JC��y�5!�����_JzA_�0Y��N�pGv�_���^���I㠏�"{I�(���(�k�o�����0� w:���r`�ML�-��#rP�NR���^�|8$#�dAZ*��WN��N)�˱>v3�hr�8�]�6A���H��/`4��mbNba�V��cp8�!4�"]$<6_{y\ ��g�	B!�j7�n9^V��]�'�$�|�u�+Z����Oɒm�%�q��Y��h�f4�#'�	��wT��Q��qE�W+ʹ���'���m�Թ�,4�����$W Yz�YN�&�	�Ņ���k�JaQdIo���U�U�
b����lӽ��|�	��h�'�<I�+���k��uY�Y�2��7>DV#��漷J���_�"0�;�Q����|�h�^�����
�����]���tIT��k&���>�ρ��U�s�=o�5��2H3{kJ�0���i#�y�
��t�?>} �B�˴Z�T�Ƙܡ�3m�ΔNIi3��,F����4 ��7�be�Ǳ��=N��^~��ZlC0w���w���Z��U��3�
�cX�M4��&�
U'���ǆIM�U�q���H0�߳V��w%X�О����I��� t�_[2���<�D�,����+�:}��|����	9��ŏz(H�u·�3�^l�s�,,�@�[����0%��dkk(������xY���x�y״��Z�����4��������i�~����nQq���[	���/֓Iz%!��$|�Th��Â�I�Lj�%� �����
BY�z�w�l��W�4�� �)$���y�/7K����XP�ݮ������MkGq!�;$@v��6���*G��X���M&`��{�oJLz����}�l�HP�k̟�CB^�6�%�_p���c�9K�#R�/:}�X/;`�0���
��ݪ�X��HO�>w��x��
�&��C8;Z8/�&zT-ڭ�I�nL�1�Z!�����[��hr'�g�8�H%6]�D(���ZrB��"/I)���P�����M�SC���rF|��ɚ�s�lȫ4�k���,���ۨ���U��V]��󼜁h=S�W�q{��[H�Z���
W�r[�d?�0	d�-:M���b� ~�t��N�Zp��m��q�H��E��yu���H)�]fIX6�=�W{�#�Q4��ePBR�fb��Y�S�:, ��5�)�_]���8<�ʳ��[tB�ި�*ͨ��U���C.'?��f�/�2�Ac�f����:Ac��ڬ3�9N",������l���^��'�DO���F�������`���s#�	����k�"�o��s�7�C��y;��i��x��L7��GȜ�����o������J��J��KmʛISr�q�$|jO�ź�[)���s�6��!��j�K���� w�����y����\Ѐ�w��,�L��8'M?kn	^�0σؽ�%��`7������W�c:��=�5(�˰B��~E�8�4��\)�R�ʹ��������G�i���bPFԭ�K�'��9K��FTN��}^��� �a�������Y��!�a��)��dA�y�l�G,�0�M�x]ArS�Ug�``. s:�p�ܥ��+Vցd�o�J֢	[��B5��TZ:�
�B��-r7���j������(�Wr�Ď�Z}zkC&@J��/Avd��j���]
b���a&�YwJ�T�0l�GolrXZ	Tq9F+rO"}��5J��a�!�oW���p�[�h����ʡsH9/�$�Y x���$��Wk8�*TS����g�.�kx$WA��j�����LioY�qp�d��O�����]�o�S_5L�˲���D�a�G��F`�6w�߸����k������i��o�����*����o��5;�(-c�*�����Ⰷ�5?�����j$;��Un��2Il�7՚Q�TqDxh�R;�d4s]���%f�E��"��BYtdp`Y��80��M(GvΑ	{�����ꖉ&��UT,�5_�1w���MО������n�(2��X2M�F3�C�|�:c��!�؍�7�5����ٵ�U�׽Ҫ&e�}vªA���T�W*�$N5�m�ҷ�ۋ�Yh��X/	�@��,�j1��ӦO`3����Q?����HwYcri6b����=��?>���B�G��W�ۊ�@s��@�@��3V��c��&�
�M�ѓ���l���0��(�i��W(�HK�:c&a��-�wEp�\r�<Q M���NC�޿� �<�u��|���1aSHju�]�e8�Ѕ��ʕDˍ��`}WM�~W���������v�	ѿ����)s�T�6�v�$��y�{�c��V:����nԐ�;{��$��[5݀I:�@����peL8��IT���*:�*��>L��~uTB��+�����D?�<j���
�Foof�/
}�w�7U�����n��L�N'����-�<�;�l�1�ܝ=K]3'Yc���! 7&���5���}����~T�/�g�;�WK��:���n9̀eV�DO��+w4)l-o���\a��g��ï�=9�?��?}}���+���W�@}X�a$�v��:V[!-b i�U���J��_������h9�]5(Q������5?t\��V�'��	�n��F١�d�"�O��x��� e�ow�V_��ԉ��T-ax%���|Izb-z�2��wq��T_3au�� �},C$�l��KC;v���%�1���;ǾPRc�,)��֓�U��u��ڶ�@9�b�*��q�-��u�?U����)��[��m���*���luf�b��W*�B��p{]w!����j��Rl=�#77(��Ɍ��h.}zr���}��DnJ�>Aǿ�I	�������~�Q���-����/�z�0���6�I(�N��
"�D��G�%��ߔ�������&����#9�64o��$i�cr%��HؼLM6�#�c��Ô&��&�lQ���ƿ][���6���Bn����?������u��c2��X�*�P��\��.�ܰ�<�c��v�`O啡���ժχ���<V#W�x�N�!/%
.�i�h�߇8ЉJ�e���"�*p�a����8�� U�R}m_v��И�E&W�o��|�S��sr�/U�Ɏ�`�>�\T���,��^,v�N u�E�]��Pl"�Ah� 9M'¬����X�:���3�����\�Xa%K��G|��7���÷o$F���%���i��Eڇ������ŽF���z3�w�@l�E&E�����I���	�`;A�$����-p'ZT�m�9
>����X��_�y3���1&�1���s��5�
�w��b�n�M:"Q2ɲW�r��>��L6�̑=�x����Nc��/W��½�~S��Y�_���e���9L��+q���}B����K���V�Q���H��N����~�I_��w��au�7�-��}_���N���RѰw��[ik���o%7��=��f�Z��2}q��xR���Jf�!W��=$��f'j��(��݃��Y�y�g�t�L(ƴq�;�C��<�hXZ���m��3[��Jx��Ux~�`m��$�֊_5z������*�Z��,|�/�G^Q&��{`K��Ðn���'<_�&�5��Y�VB)�qUL��GFsGw6>����W�dQ�򍚽E�n�AG^K
��U�Pr�+bRclΌ5J����!O��D�:j��~ v�N��}� pBH��ֵ	���a�H��J��豲�������qv��O��]����"3��l�_���*Q��o%���E `�-�i͐��ѳe��25_��mJk��-�8�z��O�B��%��JB}�<�	k�3dJ��yw�I��C�}jC+�4�/XG�vcm��xJ .�.9��6t��E�|�$!9����UW�;�ܸ4K[�n��67�91�{?�ß��ץ؏t��1���k� gP����� �_��rbA�$��.7�I#��}nҔMՠBi&&�ƪR��T�Q��b��eZ�� �X�X����VC�e��U��9F�8�PP��z��֥s)$�A��g�qVVo��9Z7��O� 
P��\�k��|��f�����ԡoߝ�;paJ��w�>����]�G-ς�E�����{,������S�R�����	i����ݣΠź%�t��\a�+F�������QW�
5���6�X�	����s�����y�nU� BO3�B�Uޔ+3�O�9,���Nh�3�\Z��K�>ڏ$�q���A�Dl���U1���v~�}c�˭�2��14�k^w_q�J��
��ԓטbXʔ�� hq+E]����a30�W��<o岒У++oّylݞ��������q�S��K�X �np
ńG>(���!�THr ��;q<VFl���96"�~����b�2������v���o1��B^��n�]&��E˖Z�j3���Y�)�
q~���pj�`w��}�X%ǔ�:�q�de����H���
���@��)��B���{z�����I5�n�F�(�e��,V���"�x��.ݘݣ��PI��c0δu�s�ύ>)S�g"-6a�õi?�1������>U3�5�k�E�ғ
>�.Z���_Cp�a?�]Ti�X��Q����|*�{V���1�ԵMі*Lu�l8�m[�TU�r<�&Z"B��a[]R^|g7�P8���ގ+��1%���;�L#�{d�A!O�̵�jj끸��i{�Y�`-"�V�� a�N
G�Xb<$�LLVݥ��q��=墅ؖv�OY�j�1|���4NZ8�o۸Q�����|��_��{�Q�V|����o�����K[7yG�F9]Ջ�W�������"S�|�d����H`�jg�}�Tt�i5�F�� v� Tc��;���3`JA�
�.�7g�D�N�Ϟ�?"�bx��UM�����&��ǀy�R��6]��t�r�e'u֬�g���Do�_�x*�E���TvQa�3D=w����8=�V�>���_�۝�JJwՎM;:'x�)����fd^���u�o1ŨB�*�l$��������8�,� ��墨��Y�ZGL�����&�BCw*U)����,��}>7�-Ǩ�4)\|;`.��ض�q���MHP6'�.�І��#���>��ͤ`�����j�n�P���Ә�v�(�a�����	+2������r��A'�d�ۉ��?��җ�^-c�/�-*j�?&�^5��!z��<�� �Sx�l��~�F)Y��d��z�G��}
����9�D.c�}b��a�v�?.�`�!����]��Ĉ���Sq�?�pd7�ʏp&���E�c�������iV"K���LTi3I��y��5I֗�q��]E�Vn�~&n�s�D:��6k�XZS��� �����6� �_�Z�����gZZ(-R���\e?�!�(����*>���I�� x� Z'բj�.Q(�zf��#���$e�L�r��r���{ǷS��� G����ɆR_q�2���i+P?E���q��,Q/w�FX��hq+��"�� j%�U�1	i`��b-���i�%lfGbQ��M�zxˣ�g@ڪ\��s��7.L����L�n��7�y�8�`pU��	�ޯ2o���1~�ZE'�$�	�)Al�Q�0�����94'#��~��1A%z��׼h��A7�BJ~z��h�g�0������s���2��W�t�Y�K��Q�M�rS�ʓv/E읩��m��+��L��+�-$4M�e
) @0�(>ym!6�d���LΒ�9�����-_�֋i��ڣ�J�=N��l���8���{&�QV�Y��J(?h�@���CR�."�p`�*��&P��Zƈ�?�}E��Y�ki�2ϝѸ_�F7T�y[L�X���e��R;������Ȉ~"�cʴ�<�~Q�^�Ǥ|4���l�љ���	�l����8���ԫ�c��ޛ=JD��OH$T���-
� k� o�Wp����Z��	Fe�'��,�0�V��ZO.�Q�)7��ph�1��R���-Z`���gz�P�}0���>*�t1f�#���b�i�\�Ma�_����d�# �J�?餖��9h/�em��K�}�i�;�v���W��Щ_�jZ�����"ڈjW�k���d���T�?}�Qu1|�j`�Q<Қ;�y4�*�S�X�!��$ek-�n����B���C�����Mp��d&�2X�?�����ur=�����ǭʒU��K���H��XS6�����U��x���c�!��"�*PȐ�a"��F���l���w�8QDdB������(�B��9hfFp��^�5Z�tƢU������3�`��Cj����u��d��[@~��"�נ���n��7��	��V�s�=D��H���o�}�5VK���DC�v6?'�ե%C��+�M8}���T����Q�G��!p�*4�h����5�W��aRٝ���&y��縋�(�Ͽ���$ʎn��^S65}��-j=�O�ߌ����_��j�F�6՘�HzYx|�%�dw[6�YA��zo���qB��ڪ��A�h��v�bb��yp��*���iv�����Z0I���~�%���ч禲r�!�-m���"�i�\ ���x�}O�?t(� ��(dF�sB᪯���{uޠ��;57� +��T��B�#��OY�\���>�Y��l���"cО�+?9
6�[<�Ē�7_C�Qo�E�3����+����t�K�Q��7H��!���/����7����UEJ�C���z�ҥļ�y@޽[�Q����M9���W'0�EG�E�Z��z�"�0W�H��}��Ws���x@�Uc�-T��ζ�jK���:� !#S�'�N����,��Kv�.U٘7�O2=U_�.����-�'�S5OX�?q��n�'��2��%.
�J��*V.v��]܄�=+�XF1n��HZZYJ3tfX����7�1Z�G4߷���DXO��Mhc� ���^AG�./j���=��\�*����ݬ��m�
�W�����A�b�^�rtGF���|j��}g6�PPϓ�joF޾��k)%�u-];M	���~N�o�9��:���V�m������<6��_�Q��[���?���r�]�2"�� p����:�a�c��ъ�6e��^�uy�#eg�cudիd�u�T�]���T�%�=჆��,ݪ(�� `,>kw����t�ԛԻ�Δ~CX|sNDe6o[/�Cm�s�xOlpq�bC�%żA�SiUڃ\X�$�P��5��#9Y�ٛn8��!���N��՜����ɷY����e�t������򂈥����;N\8jL��y��|7m@C��4���%�dJ�p���V-�V����6߻;����
���H��e*\��JZL��vB��O�/ .�N1"���E7����C����m�uv�a�Q�j�pg�I�6�U�Z`p43�i��O�\@���O�x�\����^�Br�'���}ם,H�6��݄����w�K�V�p���PD·��ۅ�A���뢠2�R�t��M�R1[c�li����i^y�U��,X��6t�<\���R�������&)�s~����m����Dy�T��(���I[D3U���^��������;�w��qA��������u:�/Ef�E�R�Rs:����M�)j\�oi���AZR�;�-w5#K`��|�GA�/$!�E�V+�cX�@���1�K�\�>��{ɟ��,���[Fu��	��/���F����jK�6d�Y�ٺ�|U��`�66)*qD�`�ֵ	�oV��d4u��/ ��jݵ���R�;?�5��Z���;WQie�v�	�o{�.�N2���U��F�mDN�mD�(*~5Ǵ� �D�;�m���k���i�<�B��ʝ�cik��)�ٌ��b�wO��nѿw����C�aQ�1@�!;g�A��O����SA�=�$U��O�ڞ��f&�VR�U�??���⤈Jc�W��ڵ�&��j��+�L��E!G�y��R����R�W�.ۘ�Ko_�k妶��6�LR���8:�Y�]e(!��i��X���Dh�,DHŽ6N���e�i��(���q�t�Y��v§�g�:� �|�{@�ȹ��7O���xeR�_�Q�c7��K5\E�fu_ط��|d��9�`�L�?��z �2��0R�^|Cw�@Q	w�c)[����=��*�_��=�yA������$�R�S �c��10�f��'P����P�u��6X�� ;3�o=�����V����-��!Ҹc�A�� ��f���l��1t�
���ce���q��~k���$�0=�wg��o����v��Kj�����n���w�-����7:�g�Q(��X&7������Fv�Bx�C�r��9�k��낗\�}_j�x��T�����P�H�;/Ky	�)V���Gl���+�I\בؑ�em�܉�%�i�_`H����Iz�k��+qDR/�����]�Lg0��롔�3���!��H��7�0L�+���o�Wm��wm����Ⱦo��1��X �I����\�W�Bj��6��VsCy����%���Ɨ؜�*ZmȸӔy4�Q)�M�>�_��F�z���ě�iv��-�C$���k���s���E��ol�\X����F��Xܡ$����qqY���TZ'K�	�1�$��\�4�mv`�]#���9��kB�i*s*�s
Z����ɶ����=X�$}8j���h��_={;��r(a�d�+:X񎲟K�)�"X#�>�`9c�'�[�x��ҡh��SS{�pZ\\<���Ѿb1o>�j�n}����ŵj2�#j1��J���W.*���s<�u�3��,�����������В�@��Geǖ+c�7�����]��Õ�և���Vԥ�*??�5��P�����Yuu�x �ܟ�ɓH�(�*elG�p�n�z�m��[ݗ�V0�u��Ad����3!D�L��N^B�#���j�%�]ȧ]$��Zl��M�Y��V�^�n5�����c䗣����>�Y��_@��� �O��X��Fg	)�;�t�t�嘦1��< ��s�X�X�r4O�W�U\��/i.�S4���8��x�F� kơl�4��G>��*��͞��Y��1����}�{��� _x>g�����)��nA|�	��w�o���D~���g��۩���k*░[���_��Xy��b��y�]�\��e[Y�Uō�^(ȓ�ۉ�k��塳0�J1��`>�zzմ�� ���J���� �O�5�1�r�k(��q��:J��4-�N���TR��r�3�
[�`7R��ۈC��'vJCl���X�j]�W)�Ğ��Rܚ�w��j�}���,Ўy2�	aK�=��%��Hb���[K��}I [xe��+ރI�y^�<G�m� �
�x�-�<#n"X�G�O�r�) �jy����y'_y�,�G�����;�H����E�9E8��V�����=�F�MA4"���T�F>�`ڡ}b�>�]4�%z��TSyaX�ɻ+,e���.��%���g�]�]MpUd��ɻn٥�^�S)m���?����p,�{kd��W���՘W�c�b�ХP��׆�\�^� gK3>�k��*��P#�A]���&Q�`@�s�Oa#��z�`{���^
��m\k�`��R%[�w/Oؗ㹬ŜG��egk��ʱ*c:0Ue���Y�����"��y3�:!1�y��n�]���m��)��/�����W?ye4���
�x�=�h<��Q�ڔ3~>�9�̬W�	�Y���ڱ3��V��ʓH�{t��37P�ḆĪCT8�Ay��#�ˤ	�2
��0�KJ�z=��o\�þ���`����7����늱�-~*�hN��5�3��=;���
���	򜭝{�o�C>(�̤��,eai;�.�����/�h۠���H����(�B<�J���������P��/~KV^Jo[Atpo��Zw�ȯ���yM���Ϧ����s=I��d����D_�*����k\:%������E�U�`u�1w�� $���Й�P�>k��qJ����D��%�%���-%V°�+�(���L�,�=M��Ȼ��,�q��DI�܍�#���@�p��&AL��+�Ζ���xJ��ʞ�>,��D1V�(0b*�IX
H�m,�[��*f�3�+3+�VPi���=�	"iɌ;${"r��
0H` ����h��گ�*qy)�X���g�O��D��{22�p��J3%���E{|��~��>B=�v���+?�������4f��W���gÇ����^�C���o�n�iV��.��dy�s{,R���nA"���wz���yn���}����S��Zz�vȧw�xkݒ�c�������S�8%=�N_��ĳ'��oė�d��|\蒈P�S��AA�H��x��40�}3_<��s��)!�cU0���.G��h3-�[��$��I��ѝ=����iC�_����J�o�b��T����S�1K��wV1w�w�Y�HB^&�q0�
g�.�����0]�@z~����4������K�f�6�Y�M68�/��`Oy��a�ﴐЁ��(��� �Q�w9<� 朇E������j;u�H��|��jZ��O��;I��3%|lE7��U�8�:}������-o�O��:��A)b#`s1V�*n�1��b�^[&��F�=%O�C#��WK�1���X��_Q�C\agtw�_�룢�N5���c�-\����E�H��q�h1��Ұ����Ư��oAk@YG��l�{:7K�������Kd/X�=�P�M��hQ��І��rqW��ic��%�S��uZ%��MQ��%1i�~������p�5AS;�B�Ay��b#��>m^"�W|�*±	{�x�'��}`�%��	$�g�0T	��LF�'�Y���f)l�(�gV��¼U�ѝ��*��)ޮ�Jҹ�E���M�����'��H,`�~~��z8~,-��R�NsW����s<����[yJ
�2*�[�pt���=j�B�̻Qվ�_>3|=�D�n	Y���k�jR�4�"
�h�k6Ц�F����(�[;��݈�~�60~���g��"�Wg�y�WlK.�ĥ���I���!=���/Zj�y��}x@��ƽ��ނo <7�oE:Ȳ)�������D�6�	�r�x	U�)?�(R��:2C@hRk#�p����p�ams�qK���u�W��%�R_�CSQ���M�.=w�����S��<����=��nQ>����"�g<쯰;g
�*x��W���N�<���F�V$�B_��v�Vl>��d@�!���`�@gN�!2�"���	��}� �v���q��S�;H�;�PY�̑�� �_��G�~�e�sp���Ff���n~�w�鷤)'^�p 5��1�D�M���%h4���`g�y�Nw��bU���ٶ��wt>���0�l PUO��Ew)fE	05����b�ߡ��R��oϮR���3�����QIc��/y�sJ%ks�
��m@ɮ������|��U�9:������X��I�vw�;��6��f�=�r%�T�q�e&vd0d�>G쀈r3����+�T�7ͩ���s�}��1�/�Ԫ�-��;�q�vj��V��%�a {�������	oؠ��z�95b�6�+��4��,���|�����Q��]Ea�/��m�����]�gm]��93�=e����z;��a����KKT����n���>��N=���cھ�TFS��@cr�3��zcY������e��(����-f�Ztv:�.P���oO�GP3��Vb�̒�p�#S��P�A�jO�r�/lgoMIX4��w��Yz|L{7~�^��k��Sf�b��Y�#s�>Q\�ꫜ�'�K�i�|O�h!��T����WM���,��5�[5��G��K�
[��Sջl��Caʨ��r�m�R��;7��L�(��a����vk��D&�`�59�X��.��9��RV���߶�x�胅��I�!���t�}�K\H�O� 4۳*�t�������\��M�z�Pӥ��/�hB!�o֥�ؓg�G@̮����E�����j*߱�(v����6��lQ��D�v�_��N��� ��!U��vY`�����ǲn5.�P
���<��#g�hɃ4��ַ"��2��h��߇��5ؑ�T$�> �h������m�W��2�!��ngܮ)�3��\��W^����t6y�	�Er!�ܗ��.�+��ce0+�>Y#@��t�P��| ��(ȃHl�ؘ���j��z�m6������~@�̖�qU���[=�:'<9 z�(-F��7��.�Ԥ��zH��Ma��d|��[�ܟ	��;��}sQt��c°:=�Z�p����eH*"Ɗxò��|�_�6y�3kM=�`87|*�;ͧ��P�Z"T�濵�o�Ka5�1h��.��K�u�#>yi�r>��8�NW��9_��(`�h������^�/5b����=�5�����8	���ͪ�a�s�_sQ���-F��,�%,H�H����G	{���ɜm0B(��$`��'�c��˷�����'̡���9�}�6K]bB�|6��B�1d����3S��wI��k��bO��ޭ�����k:�d�C�#-�!��J��g|Z ����:�7`3����"�p\{ގa;�=rF�+�?bM��/y�#1Nv��*b$�Z����qnl���W�3n�R��I�*�	a�1g=<���>�|of�Z=
Q$[�L��?}N\W\��	���E��q��[nNy��I�C~V�ʆ-�֋f���ynb�8W�7�r���R�0ú�cW��P��Y=ZM^A��D��x]�+叟q*��Q��KO,q������_o�q��晔�0(ڗ��Lx��;�5�'�<��c���+#IS�RjW�:!5��m�p%�k�v^�,6%Ӧ�6�8^G�Ѷ�T������M%�G�u䌉}�����P�j�Tw0�7Jަ�t�x��C���-vn�z���Y�1	?Õa�` U^k�)�2�y�|����#� Y��Q��e�&��~��"8!�Ԁ�_�e��by���!!�?�@#�NY��L��76�'���g+x��H�Vv>iÎ�e�D羅�l�?ar�������O5����(����������%�$��'=�<�PQ�+�n��)(�vC��e��g���l��6�Z�a��QNS�h,#�1:9��:�;���Z��W�Ϻ���`�N��+�Y�=�=1p��Bk��y�=�i׽����cP/�Eǭ,!B�s�b��;k���R�������J}{E*�x����s��Pظ>�T �(��x�(�{�����+��"����;7+�b�&�%1���)l�U:1�"��6�`!r�l92�~�N��b<����� ̥� Bة^��w >�2�����9����F\8��4c�^���@<<���d�8w��7�;Җ��}��`]gV����.\�1Z.��*��[�:4�_c~[�qi��u���aq���Gx:�D�;�C�6�k?V�V��3�pӰ��
�*������
O������8�V��T�]	��ԏ�]�F��ޖ�D+])nF k?LւױOhIհ�0My�Š﮿u��T�SL����!Z1�xE%	�5υ��o#~XO|O"Ntu\=�����^�DA�޺q:���~V_Z��t��$�s�w a�
-��y!4��}��fwT�^�\�4�:�ojq38êHɴ#��a������W���6 1i��/B�9���N7ț਽ʰ���-GUxw*�@lU���~�hu� ����O�Q�����Sw��Y���0I&��$t�F���4F�|�0��J���B�(JY��ö��ֶ�w�/oX�mbNuͮ�m�Hb�}f�x~4���a� G��BA`��1�:�Es�H��J:�|B$I��L�=5jgi-��OuxG�M.���h�.m�yu&����<Sڽ4@�@�;H:�����+
����g��>��z��]Mh�৹��~$��<�GҒEN7�:�.����M���r������Apprd�i���YU�'�"v��? 	bf��=������t��ZB���r�8�CH[tVf�Q��d��S.D���������.�BSx�?:7r��>��<�q��� F�8�*����b�%(�'� ?돃����q�N"B<;��=_�G1��#<A"E��t�Zh��(&+Щ�br��%i�
�˽~Yk'���+*���\�7���;��O͗QJ]�0(�B-���c˧p`�s�ʹզ@�<���8<ȯ(��;�)H�	�Ƅ��_C����&C����(1�{+L���"����]�d(�L��PrC���]/�<s�.��pl Mo��*� ��׵��,�X�K�#�%`����<���)�k�*0�vJ��%7q�=�S�3�1}�SS�%��ݷ��v��/G��V�?,�hɴ��wh�����dO�t��@P��, �!���p�}a*��;���b'P�m2W\U�g�w)� �5rv�t��!8$m)j���DgN?Τ�u�{�&�l�O�H�K��U�3(>|����LP��AbiyU��+Jw J�q�C��m�e!���+�:�Q㺴� �(B�K�M�`k��D$L�����u!�?��´�)�� ��c+�+
jpfխ<�0�S��pQ�OD��
3�iQyח�FKi�fu�+�S�I��� ��m�����Y�:��:���G �'\t���2��1���1I�* (�ꅿ&��A�B�xP��y�jip%����m��X(y�~��s�(&�dq8 e�=ԁ�$lYV�r���v1�? }��b����doاM-5"5�wߣ*�}���q�R���{�g�p�h���X������	G��F;��'�rf�˫�O�]�Lٕ�0H�^��bw~Ȝ��&�e���]�b�6��M�Y��!⌇X���:��Qd�� �	�4�/Eh�:�ǜe�[�� v��z�L}HYs��0-e��w��9:������u���~���cH��֭�lX�k7���(DS���I>�I��+��c�x�?�}W�e�Z|?U�tJ�"k˔X&�]���Q7�cKv�>9���h��&�5��L���u�J(%���Ad��?h=<~�r�R�2�I�N�`�����3t����}�T94��DӘ�xx���Q��@C��0�p�	/�,Oi���t*XΣ��U�8̂�1>oW�D�둧Ǆ��4��b�m^���`b߲+��qi}���!
?��K��(��t�4����w�ɤ�������ڷh,��(T=
 4��N?ϰ��l��!��v��rP%�g_��Q$~I������J(^{�x�铘;��w�t������m�F���Qk*v;��Uv�̿M�r�9.w���#l�Y�xNTó1?�1B�<�7y����&����Op`P�@��A͢5H��誷M>�g[���ޕ�V�I�#�ŕ�m�)��B��%4~�:�fb;U�����L�"M���PIPF���Px�5�&�L��&Ķ���ܤ���nT�����"-֞�#X��il�uڥ~JZX��/v��m`x׋�i�{ɕ,$v_5�ݸemh`���s� D!�tIi!Q�h)�zD	�&/mUD�Th�F����s8B�ͭX2l��'�V\Aπ|N��:1��qMbl�r����xs�1��Y��jų@ �%ʴ���8�A�Csg��{눭��@�ٔh(�+y���@;O�_��l��c���*#ۼ�
Knux�gZ$�hx���c���!8&@�gs3�kJ��GԆ �W1���MЪ���
CRӁ�'��$��������z�V�WM�f��76ł��`}
�������]��=$��RS�@��%��a�ƥ�KR��[���	���,`��ø��	��m�����D�
���k4�ƌ
ؠ:���P�~�@�Y�Zo較��l?�5zV����`�/ĉ�l^�3�� �X�|U���ؘ^C�/y'�P�W�!��.�Ò�fl	�OU�;U��몡1�Z�Bρ6� ��<t�ux=������|LEN���F0K��I�*6�L�����	��\��[U���	pP"�,�ਜ=.gl�/.rsG��(�#�#������灾��q����쒄n��$J��>���@�|9�d�+���D�+]��N幥.���4T{�b9eA�Q��e�x%U�W��M�P���ā��R���8m�Y%3:�a!!Q�R���J�
x��[��>'��{�>���kًr��N�y��E|60�J�Ɉ�ˍ�*��d�Ay\�
���7����@t���#3jU(o���Kp[��$a|��k�[��
.H�c�)¿�l�>���H�5�G`y���-���jM)G����7��Pc��@��Y�~m��`VE
2M�d����̓{�H2�=o���zz�s���7��(���c �gGY[E�#m.�|cN�?m�<�;��7��U�&��f�,�l�>+�+S�/�����4�)N�����Au$7�O�}�\i�_$��f�5r�9ٸ�9i�|"�-s^�(E��(�x��Q��
t��퀷��<���﬍�j�,�@|�&L#��f�����h�f�����K����Y}aƷB$��y�u���B�(a�X̔�[�O^z���[�z�[w������l?��h	��4�=��%��8����j��������P,��afe��S���m�I��q�;�H���0����>n����ܒڵ=sJNj0V��6W\/���R�
|bw�ʤ��v�K���k��\��/2�K�M��=R+��ࣁ���\�(?軶�n�ߧ�}�"g}l����k9-����=fs.�I9����ϗ�����lK�i( Yn�r�*�j�TtUN��mԅl�t���kd�Sb?<�&�.8M�
!-$3;�Q��w��)J:'%eQ�):�����O�P���K*>��sj!�L�ʙ�����,���9Iٳ��CӕJ@�5�16����6�[d���B��2!q�ɦ��d�j]�s0��r)��J��Ʉrt�$Ed�KHs�lє�-��'�u�0���D�U��`�l�Sjd��z�N��:���C�KN@tT���A����;�ME��|�r%���P��I�n���Z�/*H1/�|����t\�ޙ��L�:���=�����z�WX�|��N��5���G �+�5��WVpI'b��i�m�M���h�aN��P9j�v@P�c�}��tT������i�1�K���u��@�I�PM���W=�{A��8Pe�4��n��w\�%�}��l�LN�z�D#���TIN~�
mDqf�@�Ο�g��l��XP񅾔U���;�����H����;'�s;�`1��_TE�f,;�A�+�=1�
CU��g�N�o y0l���N���]�z�����+Y���,������D��� ����(Ӿ���#lܣ���뛠�:�L���ݐ}�>k�Sd�]����������25�� $�8�a�}w<x٤��C�\g�~Kfo�M���S��[Ar�JDGM��G��nt�٬�C����Y+t�'��f4��mr1֭�m\��HT
�i:��N=V=�O1#���ޝfr�'+GE���e�b�`�w@�s�µ�s��^����m$.�eىQu��+e���1\��^u��l��|r<gks����{��(�j�,�ٞ�=�R��7�ŷ+��/�p;4�����?':%�N~.�$�eTy�p��Όrͦ~hA=���fb���h�$p�o�j��X�%ONڠ:�?|-/)��_י$�WO4����B`$�ƣ��/��ȯ _@�p�p'��Ÿ]�X���K�r��.�V&ŏ.� ��/���x4R�w����|jrn�V���v�u�� ՏJ���S�޽�Y`0 %��ҧ9kW���&�}z��G��I�Q��{K%�����^F�Yf��>�����pj�fW}���:�8/���ޡS�n��w�{7�bq=��X_�`A��d�@�óe�o��$QJ���MV4I��i]�}��j�_�gu�e�L��5]�D̎.Gz�໤���U�����tA}Ls^�	VAI�hA � CI,UO�>�N\$�=F.E��@6*h��(�$�����K���"˓<*�<l3��ͫ\���{�B'���F�쮏��!1!���I�q%C��������++�w��9���0����{d7�{{�S� dh�DR�f� �]_����'��C��$�����mm�+=��E��@��w���{�
`�"ZXlV�)j�pS���8'QJ�ȿC(��-u���o�Km���ނԄ-��$��0t��a��͍����nSt��=w��agH������
Q�@N|	̒�\�D1n+�B��2�&��Հq���m��%��t0��\%p^z�} (	��8b��_w=t4��@ĭE\ �@�E�8�B�xs�urg_��ОOoB�GuK3,7�%Jq>;��C^���%�9�JG��tΠ�1���n�7���Vw�F�Bq�����aH���9�����Nݟ��}��`�n�6R���*e��l��Ŭ��=��Oh��Q�����Ye�*yJE�Bqc�����ֹs� n���?X�� jЛq��k�{<�� D��� !Q^)kH�ŵ�v��C~���(?!Yc��hM����eM�������3Sjl;Hg�b;mX5&w���NoL�~�
��ae����N���|��.��e��8
H�a��J$ 	h��V��_��5��t������Kת�QOt�R6�ܓ���� N��R^����άAw�:��)`��(��K*c?�@�?;�ŕP/$�2�AA'Pb����Ihݿ��q4�&�|N܉���djnJ�7ni��Q^uo�т�@��R����5������61��6+�淋��5�a[���ü5���s�#jv'|��@�����Cu9qp���v���c��� �e3�|tdR�š#O�2��V����a��.{%t�[�w��_.�\�c����7����<����8�8��v��\�eކ^)��s��>(�ӠJ����r8�řf<kD�W8��u�4m��9-����./��?0�#a���l8<n4�+=������}j��D�����`%�GA��]����Ϧ�7�����3,�L�auC����r�AO]�(5������Kj<w�ֹ"`G���[W�ܙWv���P���5�D�{����E�����y��Q��#(�C�[�_"�=q{,�>+������E	�.RS9�^O��
/Z}����6�P��"�d�닮 3c��Qo#�;_����}�/�NTa����b1��2�Bl��o��,][����Gp��K��IH,�����\�b���Äk�����0��;��@o�+���*Rh`��7�a���;ꟑ�[��r!�Ũp0���  �i��n���p%D@��U����p�e��51ɠw14D�L�)d�k"3f�F�{������m��<u�i�DZ�����#�;Kv���h_�Ţ�_�DA1�_+�8��B��)�3�¸�C��WO%��}MiK�����[��!��u&�#�ME���&)�u�NvQ4�'�}ݤܶwҽ�%�+�Fd���]yk��&Fb�5��Xb'�Ph�H��1̳˔́W�z�V�NhK����U4����=�k�#�X*���m�WD�Ҕ6�K�U�I�f>�9͝�rpC���?2%�]��������Me�YmU6��!�&�䤥�]�C����)ͩF�ۢV ���C;�-ze�2��[/.�y�����;xp��*j�xO���V�
5����.���9��}�������,s:�W�$w/<��&���M6N)���V�������8JoIY5�u��C�\ޜ�2�.7���W���� 6�"K�1��������G�۳�1�F��0�˷z���g�;8�h����N�k�G�<�@H��go�u��H5�3�}q�M�]s�9ry' 6����w|�VHO\�:�i�EAG���n*�SR��mu��E51a{��F5<}6蠖&-_��d�r3kLF`�����G^���0������#ᵄà��Wf�?�2�R�d^��0�����W�֍k����(�Q�'
�`�Ý�}yQO��6�!�,{���/�<.�b��YQ���>M޹�$#?�x��F�}|��K�r�)R���:@���:0C��w�_e6���:�^�
��D�]����Ez4����m�b ��b�5eo�D�iy�N�hH������1X��!�q�@ G!J���`�3q�B�ؿ��J;�k$"�矝 �Y;x�gr5V��"E��M缺"9���9��(���h{��2
����.c��L�`�ƴ��z.���U��$IGՍA���=��q�ji���Yܿs�D��$Pb�@{���θ9Tq��UOP> u� ���ztKk���z�dM����_�l�/N���P[?
���:sy�Z��X���'나Q�gj!�eB�[�Y�He�N����x	8��x��C�爰��� p�)�C�.��+����E�}��P�]<��p�nL"�����6&��"a��yA��1R���(>Q����+ޞ����u+LW��eWK�w�P��$0�a��9&�A�*��Y��_�6��F�yFB��\b��`��=w`p��+_��^�6$��b½��m۾{ŉ�$�@��F_��KJ���,KD�R��C\q��?P��w�zK����eI���(��`-`�ȃ��5�g�GY�p�LXGbg��<ڽ��.9 EאJ`�z�C���X�}wλ�,:����$M��⩐�{�����,�z�ײ���_�p�ְM��C�a��ҁ��)%M��:��.��@UО�β	et�PT+&�_,H���;U�X�uic۱�-�%�}�,�o��t-�[E�?n�\��Z!c@��F����!�5gl�>��u�9��`��SE��Ω�Į��$D��p8I@�G�V)������݁p%�'�,��7��w�:������*g�[���hO����L�u��?#�G��H�\�������I��x�������A�gM���{~Y!���d�X�bQ��gvl�5�s]�H��i#ς2Prz�y�-,@�8F�BcB�z^����en#�q�^ �����.��lK�_ikG�{�������Dx���/���N��9���2���[��2�ՙh�_j3˝ ��2F�:R�1�c��W��!�0y�H��|�
n���|�z+�r	�����[o)Abj�����(���ܿ�������P���Հ}0�FZp�H/���XD8��D 2IKaT�Z���.>�AWb���iK���x�Z��!���~ۻ󦰀؇/�	]�1l�������- ��&�;^�!���s����*�9|ȷ1����iH�$q��$ů��*� oK`���=� C�-#Є"��f%�U��m��Ab�h���CJ~ê2���R��0-��	B�����\Դ:~����f!�-{tJ7^a!_����M#� ��]fto� uy�T���Ŝ��kՍ���<w��oBn��(<'!_�Vu��B�O����a�OL:���o6�J��=���ܝ������;��W�@��T�����s����N���8VUl`��:�FT�(��/��l��QF�3���D]zk�9!2�Vhh����@DF ��;q�@(��|;d��dsݿ��9"�^��*%?Vd�d�Yd�&5�܊R�W9��1K��%�p�,��6^A�\��)�J�T��ΉK��g���-��;A����ƻ����q�z_5@?�Y�~t4m�䢲ʕ<��C�RV�h#��'�)�kU�?��6�F� Co�P��h.�_���^�2�d��k���/�W�Is(�d������f���9��~��JL��[��E_�v�oE:������R�e��A�f�Ag	�C���$A�K�d�\h��oE�Z"@��E���p��&^$�H��"+�x�X���V���r�E_�X Ѭ��<ˑ�D� �B�z�K;����D�u��Bז�}�t�π}�b�s�у�����N���F�"�Q9�C���"j�� `�h�2���Pc�����/�9]c-�����.�f�׵�3J�fߊ˓#���Z���7�zg.6��L��1�R{q�����R����~D�e��P#}��5�	aċ��,����=�kÑ����k����uh���K6�gKk���Tw��]��3;;M(���I��S%/7�g����T��{?9�����.���E:����i��G�5��t�L��쀖9y���0�tj-��4.�i'+\��F��q��{7�R{-�R ��8�
���@w�j?�=��9e���HC�"^�魙�y��;�QJB�b/W�.+5�7zZ���x���"�/�[��5�j�ts��4xdI��}*�Xg�P�Φ��=�5ֻ�,䇳�RǨ8�^s@S]���ǲYSTE�~���<ߔ�òԖ"
�*�R�#	�.�^�QA�	b�x�n�n����ͺ`�ޛi����ſ� �(���l�9|9$�R�+S(�/%���XcH��
G�߈��b!O����mecz>9�t��ԶY�!\�4��9����z���!��>���r/�aI�5p�����]���tꔙC\���w�k�h�b	Qv��O���7��X����^���c��+6�혯� �$�.�b~��GW�)C	$�P���Ո�-r�/"^�J��#��Km"7�*��@w�C�}�u��:h�Qb�bd��j��]8,u%g�����,e��(z72��HrpJ�A��)W�v�<̃�;a~qq/hb��/���T��c�B�1��8�t*�U�K���+��=�ZUg
3{=�����Pk���e���p��o`�W���ixV�Iz�s�y/Y�I3@�Bϑdt���+��C�{(Ku�q�1y"�|ڤ0�E2HF�hBbjH�n�э'!Nq�Ǉ[Xt������mЁ���[Ɋj����#��u�v�eI�č����ODh��kuޡ@6��*��c]�m#ߒ��!ݯ*/�i�]:�M���<�$�p�3��ƹ�⃂�F�}�H����E:a�:nPG�@|P����n�!	���yMg�C�����o(p�b��R��;k�3*��T�
��ǞN�:k׼�n�:q�,񺆇�ɱ�D� �����QHP������o�^�%�n�5~��:c�wd���)�Uħ�m���-s4������SW�1f�hހ�ԭ2���"�L*����}R�գ^+��/��ݝ#���T��X`�x�`:��Z��O��Ҡ䉱��L�I�De���&7��w|��T~�?;*s`����i�T=�H���f��d7�9e{}���S�#�.�,_L��R,���t��b[�P~]��H�y�����E�������kb�U��<��e��G}��l^���)
 WvM�k0c�vGb�f��&aO�n�5�������8>�r
��{�eT�iԱf�SV���OmX�1D>R�,��n��ށ��n��
��� ~8���q�yVM�ސJ�A~+��	v�UW9B�k�b-��av��GY���,T6Dq���8�նSO�%&��
p��6�Y3>

paG���ʧM7����9 Y����W+m_�u��W�ϰe�O�&]��*e��ԾKn��c�)�~��֣�_�p��R�"؅�I�;�%'?5�����#���Wٜ&��9�5�l5.< E��˶^-"F'�NU�ɕ��r���m���T-����N)rGi�����1�9ET�{�h:N�!
����L]�]э8%cIѰ����Bqר��Ȩ���N쒳�/섖�Y��~3��*:A������Ȋ�_���
�R��޸�\_7m���2���&m��� 4�;A�9�����l�&��J����#S��nōW/A(;ړ�و���v�l�v��w*,�?���i�x��Ʒ�Fm���+�UXxh�7g�[��ğ���C|8� ��c�E�{�kE�>��}�)ɰt��=�%1��or'���r�?�H�����<��y�n�H�b���g�o8_��it{���4��tf��?�T?a�4�Y�!�c�^�{I�;v�<woc`f>�ـ�KoڭE��yyi�v�е�K$Q��
��	ZЊ���P=!hL�����ޗ�l��pA��u(h��i\CPX����[3+�/}E�>O��y��q����'�$Q?ȁ�����r�_�	�8Z��2E�i�������dOP$;N8��W_IpY���Ζ��Ĩ�۠��!� X)K��-��#�F�g�H���;H(�D��+{�t���o�mK�P����h�������#㨦[�-��W̃[�x���6 ���~�������)ق]�Ӑ�eы�o�RH]xyn��ܬ����R��كTCV���3S�\5�?����d��цE|�z��ymb����,���1�SnC��Xc�<�y���9H�GEFxy��z�&�C��I��* H�e�yTV�vg��*TъH�*Cʤtv���~�t��f�%�L�?�Mqj�������7�.���N�� �fY^+軆�2�)��g��m�G!I<S]b��ܽs����6S��bX�|O����ޅ��C�����"���#.��a��SH| .$lr���_\GI�'�*G�����3��>caQy&f��羶!3�� ��v1�q�ct�_`�R���"��f��C0�re��$I�?�4P��}�:�[�pE���BB��Oj��u�ɟW��A�m�GN��#rt�|j
5���U��:���G���rA�K݄������n����S�A��1o����_V�fх,�w�+=�Ҷ�Vf��lh�1��g���:�1`Ue���?#B]��V
4�^�협�?]_>���� ����� ��GC��V���q7�FY�]kA6��3C7�A������D�c8&��V�W~�L���������@}y�.�ԇ����:� %,���0h��|�wP(J�_De̝iS�s��X:('�[�Dv�#&����R0�!�����~�Dյ��hD��n��@����pR�6U�2t�!������T����ͷԇ��
�p\Nc�F�$�\�h���¬"��_HG�@f��Ta(�}�^`�h�xL^��>^��ݐ,'֕X�%��-�%�)���n�L��z�|�Ԋ"9ޯ�m�av�c~�;=�35�r(��%�#^B3�9�����_0�x2\�$ǋ�|��5��")kāE����Hq][�?�{����;�B��FX�/���B�p�����}0y����b��s`&l�</�V�p.m�����5��X[��@V~B�̩���Y������DC��ԇJ8&��*�a����`�O�������J���Zq��G�O������ĉ�fy�S���0&6�O��>��3����
��۽���^P�d'��"��$�E{�K����Ϩ`Z���kkq�"R?��'���b�/�ȕ��'��]��ɠ6�|�о�n'5��s>���~$�QPZ���|��׮��4���H����;aa.HT�	��	��9G|��A�M�'��C�q�Њ�;�}�g��h�t
7��9��/����x]&��m�L>��2&%�����/�Q�T�0�s�tv��t��˅�k��{(Gʠ�;#K�	��y����ώݛ�d�
��Y[�#�.�}���@Z�Q0�Z�����	���n����r���X;�/��2��+M*:�kd�ώ/Nڴ�7�W|�毘D�Y�%�Oy$��Nlű�>R$��M��i㬰�a����9�3�� l�L���=eMtS��<!/<\�糣��±�m\�N�p��W9�Lm �&�p��>i �o���3z#��ݿ���$�X�{+RP�(%��\�����(���`Q
=��:�pF�I����zgt��}�_�m};GГ�6C��[�`��cLF#�j-�k�!�b{����1��D�{
rH������\�G�X<I��ˌ-��X}���R)]충�oQ�3��W�?�*b�[#D�k�����8hҽؐ�S$-������>ͭ�����_���w�*�?!RʁP=��%y����C{�Xtz�J�r�]�d�g�G��bA����?�Д�����+��"$aSg@��"C���5m�eP<�[48ܕ�VK���}�	~5�is	�Ǫr(0�'o�B����렐���>vc�x�ႊ���n�p������ҋ2���� h� xHV6��=;8�ӛL�BL#��H��݄�x~��(���̀E���u�1���oV�mAρ���6����X�8��S�� ��K	�㌋),����ӏ��v�_��gq(.�ʃr詆v��~H��B���c	�����9X�%�btA��ȸo�D�����Fʜ���n� 9���	�����|[��L�U�� -�b��ʱ�?�&�\6Ѱ,�qͭ��n�x�K�Z��$�T&0��"J{�0x^��&Z�em��b��f�0)���z7�G����;�w�}��j�|�B��UC�W���0�M�2v�	�/u��7$��Z��й䀲1�#e�0�H|r^F��@׆���H+:�HBV�<���x��W[n�f"8�`��e��GYD��*OA�����|��ދ�	��YDc�2�!�*���3Z�r1D�|%,�B�BK��M�����Ä��r�	�]{L&R�o{۸�m:���f�-C��H��c�DS�}4�j	;5�[�/��Kk&!�Q���9�H��]O`�]��I?<X�*G�+�O���]5svv�;�m�e�jl�D�2�P�]�)�z��+!0��dVi(�'w���PO�\ /��k�����'�k*��*J�i�e��/���}����Op=�MX�2�&Ȗ�5�ɔ�X�\� ��S��D^b��6������f̐��_��ᧇ�j�ŕp8�}���lX`�������.�8��I��8�LnwyS��Zc$ˋ4�G�������s$ �����1�̆����[��)����|��j%A�W$ˮ�C�57�e��v�I�� md$����A��P8����Z�P��aB�dx0��xbG\h��0���_B9 (= ����Sw	;��9�8%��yi�&nSK钚��@�^Y�wr�_�C���9v��tzS�Z0F�P#$o����-<����+�UWJJ�������l�Z�M��2���7�M2��h�l��ëD6A���+ߐo��8�fV����} V�ns]u����~�S7q��L���SA���5�B�,<�\��,e�[��Tv$�^^��J�v�G'�+ݐ7�N�*h���zO��S#Y^����)y��9)�Y���2J=γ�	���4�٥+����K��,�K����K$�>�
['��{S��G�&��"cPc�b#��g�}�C�V'V%�U��տ3���@��f!�X4i�IbՑ
vg�'븆����V�8a��u��p�H����u��ˬ�g[sL��ѦdH���7�@2�\M� :S -]��x��T�72Ǵ2ڼ����DH��O����o��������*7�B���~&?`��qA쾏7�])�:�X��)#�qȥ~t}�N�c#��YE3��F�F�Re�x?�s�g��Z�Y5�f�w	*t�@��	$��'����x#̷�墌m7��@�mi$aO���K�q���C.�<ϐ7B��JB����1߂�	�d)�0t&�	ے�Y�,�Z�"Ҩb�����3#���~�9��\|\�W�>ϻOH��g�(����Q�*J
�5
���V�,�\?h8�����]c����u<)���z�JXn9�w��u{aC!�Xփ�X�{�;6�)�t_�{��Aa�d�%�0�-R��|������h�f��[���$��C�"�V�w�}7B�|��lr$4���G�#�<ɣP�1l+NS��7��f�Y�L���k���$A�>.�Kt���dW*�3���]��z��I'�-���[������%�QC��(��:FI�D0��b��Y��'�!�ߌ� �oM�yP�0�`�zK�d�GI���}�􅠟�fŸ��x0�靁N`��r���HS�%� ���oǌ8F٬�B}�÷��`z�5����#�C�p(g}m��1d��=8�ץ�2�`�|��C_�,g�ݨ�������F��E�;�Ze��%�:"|�:<�*��(����gh�B�o��e��o�>��ܚ�Z2�G�Ƽ�l�$��ܭ*�L�!z]=8n�m�΢5$�,cB���U��H9)��ʕ����fEm�_���/����AR�����.��Mȸ�����a�����:�h*����9QEY��v��9�1��X�~��W,���<$G�vQbw�Y��;Px��xKf��W��0�4��px��2|>��<�A��_��6�����K��&C</��p�K1_�+��Ҿ��/K����BjzJx�o���f	�w�����n"��{�~�b֗����v]���m��L9I5v���X�z����A�~^ڊ����i��ɂ~�G�,'��Iߔ`>��BX�fp�%v��4`���Ů�%q��%�`���5��Z�{P�pjO�#���!��մƖ���8"�D]YIu��V�a�T"���W��	�93A�B�I��&^΅�=y^��޶�In_My$�q��i�J�ԝ���]�G\�K��$�~8����l��T�O �ȝ=B�qV����0�34T��˞{�;�4 ��+�|A�ʁ'��` &*��N��[ �R�h�������\�cU�h!���B�����@�\��^�E�a��0�'�̛��	��őv�3z����,� x���:�o�@7-S����/�x%��v��n��#R�Eg9�˲)�>Y_�&&#?���T�?����R@I���!X����-o!˃��z���I��m��c�ӓ%���X�l_v�������)��mb�^{�}B�x�ȂrռFa�#�C20����x�������X;�0_B�$`'�Щ��bX�i脞A�Z�6#�'�6���z���>Lݭ;
��Z���ٽB�O���%��WP�Խ��t�`rf`�H�����#�4���tk׻��͞��0`��Pϥ`^���/�v���c����H�D����DB��n
c��䫱�2ؙ�xR}��[俥��|\ ����W@MH#ҍ�վJD=�4є�6���A�'
2�Dv����!�'�#��f[H�4���z�߶Q�5�8�P�6K��1�L�Q7ľ�J ����-�t��1�Gǃ�']�"�lp��n(�^�F�ti
����((����m��1��R\l�uA��o�B=�H�Yd�|v����g�d���Z�P����S\���LiB���@��"a���s��R�� �W�)���Y�����95�!���D���7���u1�4Ͷ�*-��,��t0���
��UU��M��q�^�Nz8Oq�0�"zW���,��2o���'�%�e�QT���)\n�������0�?6�A�0|��#�zZ��6w��\��A����Y�C^G�s`khogrZ�<#)�����c�jY��\�ـZ�X\�nrN%��6�a*K�?�l�z9�|�7�`�WL�=F�cx�YI���z���'�w	��[_]pA�~_ɖ�l��0�+�����P_��*^��\�����ʿB���|�����W��@u�}�P�҅?4s~���s�����"�L���;��5��w���Z��}���hH�W�&�����o�Mz�ؚY@1��t�{5�{��U�l�CםKh�]<�\���X1��d	<�t���j��,�s�f����7=��I"8-rf#c�X��]X�M�#��'��ʕӨ���~�����;�S�i�]м-�pӐG��<!�	��7v?q��{}oO�̹�GE'S}��ny������D��'���j�v�8�)�r	������$�$�ހ�Na��`-��EK{��l�I2V��y)f����}t	��(�9�	�O�(���#	{8]A��
��cؓ��i�p(k�DY)�p��G�8����u����j��o�f��s/���s�u�m�ε�:|��t �9��7�t��*�Y��<5��Ȑ2�7A!�L���İŰ�2;��mK�o��7vɥ\�c"*{�"q������~��ر�88��()b�Q�� ��	�t\YޗD���V9�u- -'��!
�	����$z�$���]@��ˋ�k�����<#C�[�8�'k1K+�����<�D,�O���\�E���^LϷg�o�δ.���\l�>02L��"��~7�'\�ac��)5+�IB|:��3s�O~��V`{����]?ib��`��a������%�\��p���9�oy7OY �Ð}��u4���B�0�c;�-�{������'����N|Df�J��Ǭ��J�OC��I��.V�]���WF���{�k�ZJ܍9e�v�q��ɈiYC�J�}�����r�lA>��y4խ�<�ٻ Yϋ���7m5~4�	�*�h�g�}�Li��X������i�!�u�����E��c�Q�³��;���&�8�i�f5�ퟥ���~*$Z+���/*��b��Ks�@Մ�/Цy^,
_��kN���?̿w�)��N��5'ʬS�k1���j�+u��)o�ʎ0�o�I���S��DN����V�	cą���L�y��y�ػ� ����[��X����&�M�. �R��m���)~���`���b�v���L������62��Aa��lֱ�.�o?l���G�������.�䰽 !�g1w+���$ H�2�����a�v�J6:�I��gz�'�����k���o0��/vY��޸�us�:\��	Q?�C9iMo��C�u�?��|8y@l
eKJ�
5HV���4�6}I���7�5���ܯ�p��%"�ӽ�wE��〙M4%����R��S�,d��V֨'���zF�m1"�X���j?���)��pwfѻTe��7d�/�I��?d`Q�4�����G�I��]n�G�2��a|��6�-⤖Of�J�*���Ǣ�M��|�:�0pD�a�s���v�%�AG��*�~;�Fþ=F��R�;A��n��{R��f[f�n��s�5;�Q�I�M�Q듎��9E�����K"������5�4��oc��r�_���ѯ��3t��g�*ս����̇υ*��1W�o,g.×�hA]E�I�M�`꯳��+%�
o��������.��h��7�����HM�����w����m|��y����1vcc4i/���wM���&�P�*;I�����)�2���U���`�!/ư�`�3c������"H�x�y������ �	����N�>�M��Zc�-i@��r�܄s��1�:����8�f,�o&E���}->0[�	�VeӪ�
B��[�:����
����#��e5�e	f�қ+*�p;�#�}�Iy�:k/t] 	N����7
���ʭ�T�r����v��PW�t]�����A���`���
g	/5Ep2��'��'Oi��KC ��G�X�[^��4�%��O�2|+�5Μ���9�	 �Zv�|���έ�ߚ.�&��У�(��ᕣ�Z�5{ (iW���Ʀ�{A48p@�6^�{Wx��򸜸�Du�p��5?�_[O�5���:g̶q��%OAf�8	����+K�K��h|uJ����R���t���l$p��X)���y�(2ݯ��X��5ĸ92�R�A�F��D���C8
τ����I^!E�V�������Hݤ>�y��Z6��e%y�k��B�oO��>�k�.RL���Vx~8��i=(���v��Oޥ����/}��k!ɹ�K����M��X��K/��P�o�L�d�p�$B(%�#��̓�SW���`n G�d�GK}4���n���73��u��خ�;�*?��lP��(���J�#I�|�&�W�ɪNε3�_���{��m ?�OG��A�CJ #g
gӤ��
x�R08�\�����wI�s�
4��UmWۥ�NE��u�<8@�JF�]�X2��/t7-=�����/���,3;�D�-�l��!)���tj>y�;�-Z��8OdZZ>�Dy�z�K�}6���Ko||��X18_[K�X�%����ʑ!�ٙ���l���t���T{��C1a�y�μi�:>�a0�^���s٫�>#��V/?pm�������p�6_Y&���/R�V��n�ޙ�������p��Y������� g�p041YmI��k �����K�K�6�r�I)�rs�{�*ڐq$�s�A��i�?��rh(�	m���p\sg)�6
�*�zG�>:G��k䲂J �LjXއ�+����+M���<�ulp���ƕ��ޫ���D*~�;5�� ���!
�S*봺h��а�
hb��z�Po��aM6���w֖�	#̙��s��:��k���?].���ls|�4����}��6̀~L�/Rc��&�JFG��'Ǭ$�Z,���	HUď)�x�K��u��P����o`)���+Q�+-̈Z�.bmC-�F:��0�
�}Vn�=+&k�tw[�+wD��wXp�lwq��C������< �8��h�]��&��h&��D��a���Fo+��:'wA�6��@��^�J��滛����Յ�Ϣe�s��l��3����n��xJ"�G�p��B��Џ��]��
 ��@����eqB^SC�y]ә��+B�>n>m-t�*�X�7��@F�"��JϿ��x�����:>�Z1g��W{��a"�I��X�Ч��X%��1�����C����œo��	#Zi�3z)����f���Ƹ����&�S��2D�KK)��ݬՃ	D%�I$^��:�l@��J�}�Di�T�(����.���ѡ�G�΃���4y���g�w�"l�(�������'rq:�	q�h��`EI<��wӅ��a�����p��\�FQD�/���_�Y�����dq�s�Υp����N���|}��/�W��E��~Z��RB���=����?���#	��+��Y��n֍ٟ8"�ּ/M�� P�'�\��{�[_?��ƢD���y @փy@�ݚϷ��lQ�Ҁ��Z�m�V��E�9*��)|y�I�J�B�{��w��v#uҷ����	���W �Ҽg��Z%�����4�W��V�^�@��^��_��W�bF�@�Y;7[,�^��dc�����-���ծ��$�h7�wAAj�J���߆1�F���}c`C�>��M��-��\�"�O�F�%m�T��h!4ǌ���(����=����ʞ�+�b�AILB6�D��q��:8��È���.�(�X�`�z�)�"�ו���)ȣ}�Td�E>��y	5�&1c���wE���[jz����O�p�h���7�����z��Ů����E�j!h[1��VB��@a1��PlE6;����(_�3�](�:)2�Zj-����ls�e�#��	�wb�-��]j��&���ߍsl�x�ǀf^���[��A$���Y��>��Xb�ךIdWץ�^}@�*���{A	�T��l"F�=�����>�EKU�-���cYoA��5�0һv���C'�b�Z����+���;J����uG��{9�W���T��	УaI�ʠ�lf3������8��?,Ev�EG-;eY��qgL��	��Aa;��Ǵ�f�7 �yB�9zbe5F�t_প�l(��~N��{26P�[�|�*��ƌ��	+�~�PK�le�r5("���>���=%*6tW�ץW�U+ _�òB�� ��^�/no��5�k�O��o.�� 
�2^��3Y	���{������q��1���S F����~��sQ�]����Z�p���GV�W��{OݍQ^���[͹��CO�����a�3ų��l�@qZ]δ���}�?��5�;k��7�
�)n�KmhA���Vu@�����E���)T"�r33�ܩ�Pm+*�8��b��aXq�,
Y�Rf�pj]���/��R��gt*��ګ;�q�,1
��+y5��p��%��)蟟���-�?R�)9/�F_j0��z&�dG ��L<?��ynL?�Tj��;M��fe�ZSS��b��F.���.�W������R�ې_�!�d�v�5I�w4 ���B�=�w����������1��33�k��dff'��-��=_���#�/.-�|�ơ4`?Zo}V�]H��6���4�WMH�aŗ+�u�\���E���*/���P�>ɢ�e;�k �x�֛��P�"-5ޖ� �f���r&�xg�����E���&Kt6�KvV"��J_F
����$S��n2���-dv/�eHP�D$�u�J�T0�/j�5�]=�Ul�. �FB]ى\�5�>�^I^67�}�~#G~7]M ����?�1�lY��;�&�9��D�8���?Lq���?=�8}����}W�������AT�iQ�n�5}u=
��ܢ�t��|�fr`N��,���rU��
��a��&�|�Z>B����c't�Q������ְ�{)c���[-�vǽ������+��ē���ѥ���4kl��S���a(������f���`;���S���ݖ#�Y��V�y���G����۸�%cw��L�H*�v�qk�'�Z)�n	͕GP�f*�p���;n�j>Z?zbU֢^[kr>c���;�������� �phtYKUR�*��$_�r�R�֚R3X@�"���N)��^R��t��)�J*��2#=K�ʚ裱��"Z��W�r<�A����$0�����n��t��M�.��Sw1e\Npe%��ೱV�{��*�n�� 0:��A�����|��#b�ZO�Z9��A\��>^|' 2B��n��*�FR���!N��A&�m��JVS��&����=��{�Ԑ#q*Y�������C]�0�tnva�v��bX�;���9��#j3��QlWƋ$3�x�;��M���!5�C"0g��������p�|���(��N���͖O��-�}%��E����K�ؽU��'�Δ����3긊�U{�$�ʳYmɚO	)d���_˞L�v��]��@}�yJ���D�� ��R4���2�"<{��d�C�!����6��J����8� ��,i�9ʡ��@���+�` ����l�!�&&	�dJ,k�����4���T����MO�f�!�P��Z��#F���%�|�f���B�G�4"!�v5­hV*v`�<ؚә����+�N���O�*�3|W�0�w:Ծ�׺���%z�(
��tbnKO���z�<5ݽ^{Oyl�7��N��O�GJz=�698�O�dV��8����T�!�A��@'TX7Į�w��<4GW-+�VG�6�����	խr�x�ޭ�D�W�γI�$��`�͸�ݷ�d�@G�bʳH1w"�����h�>�c^ o��}x��#�`�=��(VS�Z� ��*Ja�J֡{q����.���NX�v�U?���Zuc-�`t7�*��@��)-tq�C�5Hr2�DFt�mW��g��#�%�wW����AR燦E�^�(ָ9������%�{��I�Sօ_Ac�ua/"�����g���jŤX�d����X��땧,��
�7q�����KH8�؛�R�na�9`<>�z�P|�,=/2`}�d�}ݰY�0���[ �����J0����_���ć�A�M��]>�������ߎ���r��9Pyi�|�9�h���8�'+*�,�yc��f���7
����'�|$;�0�O�.9WM�AXl��<S=\S@6r���c8~ۢRG@�����	�o���u�;���:]��~M���e�⻫�����B��v����)\P����1�Z�>�ˋ"Z�2�CR�,� ���'h�\�A,a��A�6n`�� 0�����������ٜN��}�4����D#hN�1u%L2�B%��Y�n7�����\N���6��rpà�$����9�3��7�M+�NS��rDIf5�>I>v�!�R�����ӧ�?JhӆVE	I�\ W�G)qk�Q��
A��(��[I���4؄�u�|��]�}���x�E�'o��� ��O3�C��ť��o>��l�������Be��:���2�Q��	��Ɵ�	1�a�Ԣ�_�k����j��;K��V���{^q�����r;V�/h��(xE��c�ո��kg�YͪA��؎�>J���ET�;8y��"�B�I?l�v�r�	�� �X�G]\��������X�����'��\��4![�E�<Y~Ǩ4��P_�oK�o�Ø���vvS�d�� ���Ĕ^~��حmҜ��7��k�h!Ւ�/�p��s���Xi���f�9Q�$&
ǚT-����x��%�E�/����sy�Q�p�˯�1�W�ܤ揓RB������-KUXlG��v���%#w��I?f�ώ��ќgXq�Y��C�+�u �m�'mAG�xPM�ô�j�_��z�����G�J���/� _$������J�Uz��\.*$�;vv�{������|2��1�7g(7���t����_\��}�h�S�i�<�I)"��_�t�rP�غ`\��)�B� ԭ�P|ȡw���&�ud�a�J�}��e��I�J���1�������Eδ��d�N��p�S\�h����ؠ�iN���F)�ԕT�x���rUFM�������fa�&��F��_�7�h�	�C��h3����}�*	�K���t�<�润�U�����,�Y'����g�rz�j�'��fH�YpX�9�zl�K0:���Kٺ�=���?di�z�9�U�"�=�5Mҭ�d{,bȂ��}^��톪�|�С��b��{�w���$�6�]T�ň�}K�U����)B/S���O����R�8�,�BQԂ��JZ��0�|/(�B��cqQ�J�4��t�[�Lh)�6�q�1}��"�]��f�#���8�KO��8Gx4�C�D�p��w
���L����>��;D}b�_Í3<�Ƃ��Z+�����YX48Y�$��y�>�iaa:3�9!�b�Z��I?�2�n���Z�/��8�N�j�g
����ת�"��K��׎�iG���S�{s;G�Ъ_]�����&ϫN�	[��nXǇ'�w�a�E��(��[��A�tt�Q��ϸ�5_sU���͌N䶺�ʔM��C�.z�g(w��{}�f̵ؙ��F�j\w)��=�"#���*H�4m���0�RB}U1BMsb����[�/�gK���恷4\"�G�9
�^i��n�zy�y)�AR:��+�H��s���R�Ez�\��g���1�`/�Z�����ʙ��ifj!	+���q.�2�j��@ڧI�-=DԒ#��O���ݙa�*wHy�p^�ɰp(��a���t,sG�Q�;몣HR��`܎����2PH􇖳���}�]`5
�\�YM61�*��)��A:����&�ch�b�@epw��.��`��`���bL3���jDt� ��{oj|�C���<�
�}2�$�;R��ԃ˚�kq���Q9�jT����D�8��I�:�u=�6�|
B�����c[�NT��M�e)������.��)4��&#"��C�L�~�S�X����U��[�����!0N��Z�̢=����qx�T?_	��Rm��.u1��t,�^�`_�]������s�,Y�CG~�e��+3&#1��!�����
��w�9�d���N`o��?]݈�Hi��L�E�IY8��*u0.H��\���[�k{�L`��/�F�����o�D��+3e��e�T��|�ZBw鷓7�����i2g��&�m�y5%c��s�H�r��u�����{�xf��iC3�#sq����Aن1��w܊V��t��[�%�e��ǃ��>zp��T9������ޒ�5�~_A5���oQ7���:YZ����6�����Sw����IUr���}Lrf0���!��&ʋ��9,-�;GrJ�c�2���`cdD �������t�R���l�k�`��b�-e���K尼q�K�:9���I>�����O�N �.�Y$���sMjvxg��NQ�!��\f��X-sI$��7�i�>༱�8�D��"*���ح#F�#�rɇ#|��\h�[K*��c�i �����R�N6��I���U|w ��эP>v��p2�&4f����w�k|Pv�Fx�p��_7.��v�t %g~ͅ~�0{�1�w���? �<��.<�bz�AH�߮{R��?6b�cX2:S]T��B�:=�q��T����]���b�u��f�5oSCY2�+�cB
�M��&��m�v�]�&�\���<�*��MD6Ղx̼<[� ���n��7�^=?�<V�������C-��&���������a)���̯㲵�=�֝y]%əj_��y ;ڟTeZ%��}���A�F�ʈE��"�:��^�C-x��3V�}�j�.�&����Wf��p~���P�5dS{|{"IXZ�k�J;�Q��$�{L�4�H�,���"��0�A�b`�:ݵ���6���ȇ|W(W�g�%���%é��-쓀w�+`�ٷ�;���R���f��KO7�}#Q�E3�?��Ԩ�*��L�$w\6%�y���|}V�4���Ǳ�_x2��p=e��TW9qOpw�^��<�P�!�M_6�	=ៈ�?���ͨ@؟�DPKv�V�8��Q��
�L&C=[��J�	E�X@�[W����ɇ�Q�*�������SHR��>�U�`�:]z��! ��KI$��Ьy1 ����J�'5��j�RD�π�cq��tT���n���_e��{Ċ��=9Df�P�8�?�ʎ���Mst���[� �u^pz;P�R�C ��ơ�Qy��`���?�5��ee�,����hg֔J
Av*1��0g�J�����8dH�뚭�˽�L�*��b����+(�N��٨�m&�J�����͢i�؝��qf����$l���ۼ87tK� ��,b
d�I`"�L�ȴql"�ϲzp5�o�jyj��<�ܳ���ju�rP��O�?E�G ����ިR`����d$e0s�{bѳ;"(��l����6a�CC(�������]��?+ ��g��Mg�DFR�|�N*�����t����U	I��x�2÷��\��f��A�=��ה户ȯIVP}�(s9��Qb���a���v#2Q��n��LR{��ʅ�T/(Q�S��M�
�r��-�\����Bu��kqQߐ�Y\�ogB�#+he�����B�dv�Q�ɕ��E�������gl�o�C�U<��g�,u�0����$��۷���Gz�w����2�܌s���'������-�����������s�F~�~!�D��0���f��z�T�W���Q���Q֛�̬�԰��Nm��>n�I`���\�9i��{�: b�tѧ�˧��Ad?"��g��f����8	Q~�T���d�j���=���@X��zJ��������@�K��1�(���l"��m��p�������F�A^�v�8�y��Ct�DbNR�ы
��~����cj#���}����H�k���$�#
��b=��Z���?3Mv谕����7Qc[D���J�R���2Н��/r�˱}ۆX��b�_ ���D�=��/\�f��D�Xf�	���} ;x6� ٌ����OJ8#�=V�����i�Y����\Rn"����f5��f���>�����1f�NM�
]ן�;c$�.�
^-����!8m��s�8C���2�"�m�խOU������R��Q�~�	�������Y�U��@�hi�-��,� ��G�X����阓xz���$Pz��S��Sٕh�;ؾ<���~n�͸ʍ+y@�z�h�'�&-m�lkR��&�t�y�@���Y�v�/����:b�\)y�Ȫ|�G$@v���)�[f#1G3πToE6�]�@/����v4>\���E�Z�7W���@�_��i���؆-
�Xi�@�ua�yruR#�ނl�{���U�K;���}�٤-)�P�އ2gϡ��&���3�K�@BG���X��9
<����L8��'�4�F�����H�6鴧��b���Y�z��	7�8|�|��أmD�U��1s[��"�v���	a���^�j��eL�R~G�>I_�H��td�T�ȵ��>Q�)Y�p܁���^]8L"tRW��pJ0@0�$�<�{���,��v�@+�cT�'١�s���k��9�ዠE�]�
O�bq@~����.P��:z�M���G��Ir[�~O�dc]��׍�f��	����`rxc&"�]�K>�7�����B�@$�?yj6,�wͶ%�IJe��X��i��(]xH��P������j��p�@EQt�頃�����z����P�����U�3���:3�v�a����W��X8qL������f�X�%�ܧAP�=������t�_���
��Il��e�SB�Q�
��T�ɨ b�[�7sW�b�;iܡ�O���_¤����%�EZ�4!b~����g���7���'
}e�i۞��e�_|��#��@�u���Q_��Ƌ��*��PMk�2��d��\��
W��ޤ��!ơ�z�JL,����� �����]�|�P]�0&�m�c�7c}U�Z��M؉�&�^�$�δ�Q3�P�3��f���� 1��n3��ոi�ߡ���H�|��Z�u�o�H����\�F[�/Hs�	��H~��nveh�j�fY��#Y8)��/�himDSh6��DG���Ƀ�(d�)�y�4��*�� 'a�sxq�^��%L�q�R�흅%�
zړ��?{~��ӟ�*n��y���S�ݬ�<+2��âF	����p�x9�<G���C��]e��j7����c����iN%8���@���pxhT�epYW6aR�s��]��e����= ���w	,
�a^����0��;oj!�y�iŦb|�XC��E��l�P���+�u����
�D���0O*�ø�>A/1�-1�mo���<N�Zp�&�{G�úIl�qI&�֘ۛ��Y|�W�]�՗&�iᛛ1��'��kj�55ZՕ�Q���������^�y�Y}��P�&�W*"&]!���6�ఽǮ���D:CH��a�@NP47�c�<�f
�@�#	N�A　�/˜d�=���K
#Xޒh��W4ۉ�%2��O����'�;2�KU@�g�4�
��_5�hl���T?����h>�@����&���[p2nd�[Q�f�!_R�;���\�����*6�g*R�2G��|��Xʻ��H]Pe��,���ҥ�86 -��F!R�)fU��,��fF��#K@r�'��7�������垕�3=c�P��0��l���c����ݩ��J��wr�[�).�k�R:{lK+	�7i�g5Ko�Rs9��������mi�'�(ˆoH,� ��xÛ�n:�.D��/dw,o�'�#T�%�,N��T����P�1Q��e~�0����q���q��Z"xN��K^\@��m�E��@�MW��̆\_����P�r�Y|C�[oK�?�!ԩ�꼂��WL�������e%������Fiʹ�Г�4d�	x�@iJJ&[�
,wm|���K�@�E��z��MP��`2��I͇8�T�5A�i�&�&�8Wbo�CX�4���5F�],"ܯ�G	��tX� Y�Ԩ"$=g~|�G����v������$�&;{/w�]YU�9�R�f�}����}ǻ�bl����1{GG�U�y�a�2޵힯vP�
��2��}��� jz㛶�{(1,�0����0��#S�T��Z2�O���(�����Jh'r��1�_�aNF�% H��,hx��5�m��D��2�PUs�b� weA,C�M
������cF�!]U�Z�dF1;������kg��_k@�ƺPʫ��%�\�D	Q"t:y�2NBy��GB�>ԍ�W&��hy-dy�)¥��\J�θ�-�1���X�� ��>�[p0C55-y
D2Y=�!A�!�|����A�QV+hۀ����im��'�� �>A��u���Dw*�w���yL�<xw!�M�1�c{�?w��X��Q��[�e �3�<Ϋ"A��N����S�.��˸7�>UѴ+�R���VF�Wv����~"���ě�>��I�����d��` 28j\N�P���Lpހ��ʯ���k�A�6�f�FJ࿼�NRh��,�h;���@!
 9����D��芅Gc��?t�T�JJ�8�b�B7?g�XqA�~Z"��L�� �{�ѮL>닠N�[�s��x����^eV��D}LS?��x߫���t��l9�{tx�G7�G5��I*N���ЈF�̗�Ƒ�CY��þ�N�=��׾v�A�՛m���'�O����L<�/.\��ub����l����)S�#�%�jT�O�yݛ,���e�G��moPm aT(��֔��6U��e���ӑ����Z|(�=�q%Au�͘�	��/�O�����K+<��W_e('h�.�fIS�3q�G>��s�;�x���-�O����sG�Ql)|-�0��SL��`��W��7�f�b�C�S�m���jme�Ly��\#�y� 2�@���_�uG���b���Uep��b{ϪꔋD*m�ڰ���6��X�7��:�B+�J�y�[C̿3����\;�i�q���tu��"�u�Fv��%ӵd���c<�;�f	�u�$Q̇格O+ɑ9Z������mz����+N�~n탔yS�����H��i2��rk#������~I��	sc{9l�޿M��Fw�tE}�$X��L���x�W�g�n�r![����|��2Y��g����?��ϟAMP�#5OWS�fY��S�>���BY	��V�%�[؋6�7���X���4�T�����F
֪�imI_Pxq�~���`+�7-/�~�tV	������k")rO ��P�©=���+i�7zo�ƶO��2��:��ֱ3&�IP?�)�:�.�
h�0�V	�Y���Xt��v�X��o�q�V�1��=Fp�D��i��4���s�$�!��ϐ����ݕW8c�1HH]��ϥ�l4����,:��4�?��p��0��7Z~9������<���$m{0f�������cg���$��-4��-ꔺ\�Oy%�TC+	��Ӫ����J/(��T"�you�Vc�¬x�\��(����]P�z�"�7"��t�n2jdO�'����?LV�i�]m,^���i%�R��P�n�2���QM��uM��U�cvr@Q^�7(��V���&~��#�<�%d���1ڛ�|$V�I�Ӷ�h,�����;|a2Y����`�㮎W1�������3�#މ�B�B�&ٮ޻C�u����USi�XG�=�����)z��0�fXl���k`�9���5����SG5h^�zۊ�k��]����N�`�i �W6{c	��Z��8It�-���';u0�#*3xL4��2�'�����$뱞��XH]2&XbCh�'�W.>�+��S)��,�j�6*0!Au/��H/�<ƨr� wU�οL��GX�q]�n��I�ࢭ����fϬ5/�|���_4��`U�I�H(�{�N�a��<�'��N2�Ua�m�6�n�^�E�;C�qК��jgh�)��xkLp�#���}M	I���,�R8|��'��И0t�����LYF�����_������E\��\NB0�!������o���U�s�9F�o�$N>߁�V*�Y{Y�{xgf��8|�e9�5w�[�j��+i���Zw� �0�Dxt~ �@�sZ�D(-����w� ��>���bȪ�;������B��8-�h�IO��������\ 
�J�T�A�kldn��4�3/��8�ʖդ�%�1hUJ���0��ũEl72<��H(�4���@��1�p ��Z��FB��8;�����[$`�ƞ��^��i�w�Ԏ����I[ki#��պ�H�e�Th�	�)!Z�4�r</�d���$1��k��e����������v���R,���A�;}JΝF�!nkѤ�q)O;4�CMBO�k�	5-�Ώs!�u	 �{��M#��E��~�}P}_�[��.�{E��͚?�R�'v�5�Ƙ��
�!�7�2MW&!wH."M�}�r����(�Q�s@ �H��+�~J��i�>��W[���'��ʨ]D����62F��LQ/DYg!7�#�;��dα�(�`�����:�g4��R��l����x�K�Fj��m�-�ٞry���6�I���~6���lE����C�?��DWM$��a�|#s�
1�e?��\CA��S�[���YD� *@���i�eQ;`�[�oB�p�3�A���Zk��K��,��$��6�VJ��.�7�ov��k�p�ȧ~�e,F�6��V!E��)7�#&�ꈃ�(�!��$�!�z�r됿Ě��@�BS�`��qC�MK,A٦�j��լ�2�f�8 �klP�����$�g]g����dl�e�s���$m�D����D�X���Z�� P2m�W�~9l��{����w��qbhG9sX�b���4��6l� 0X�
����������Ɛ{w�N�k�l�u��v�!�yd�!��8t�Сy����a�l���h�]��(;�SH���#�\����ݓh.鹦R<����`�L뜤D��|f�$-s/a���u�uΪ�vm�vצ �<�Ԋd�{�>�I�[A9�?Ns_�v�o�h�y���Q�E"��wd'R�����Oʹ�	�b�i̩J:uN��gF[p?�{gy�� �Ir�|IN�l-��W�_C�`N!uP"2�Y��.	�i>˖�.:�/>��~(9�.)��ڬW>(ͰU����>�1��k_ꌞ�����[8M>w��9h��{�c�	�y��݂᪞���٩�rB���Y`O!�ŋ��Z2����u�.�65�Րm�iX��U�I��*@(���(���%�!Ғ_l�oE���U�I���B<���a��<3tT���1Ǩ%�p�T*�}��	i!�.T/�&1gI��"d	1��9 ���:�J)�T=��"���D� �$-4���+�ZK��5!��m6�Xs�k��W�Ki0�Q��!؀K^W 4m p-y:�J�ܧ�U!@��lYlb��x��@�_���L�eF�@�J�)��T�s?@���t�w��{�K��9Y��9�+nb�&<�'A�sB�(�ƙl�׊0�����7�����g��2�Y��ח���I��n��w��U=��DgR�ԈE;3��8}��?��2ւ�$1��5��T#�$pҶ ��ݰ�*c'��a�f\�ʔX����i5S���iG�A��~������~�Uѐ­9��/���F�(�B�� ���ym�m6q�I�$�Z���V��~�������Y21�F�MS�u�V#H�UE���@�U�}N�5!�i�W�߳���?�U)��y|f./��4�@��h��"�-��'X�u����#<R��|v�/Z�ɬ��wU��F���@8�C��^|�*6]�D�}Y^��ж!>͢���͗:(����<��͏��5�%\@ ��#YH��E��}��_���ϻ[��Yb�+'G�Ǳ>����9�������ڴ�4�*[�i񴂰��"���]z��4��Wo�P�,
S"��J?�/���|������J����oo��F=fx�u�m4<3��	�^R��p2)R�;p�%_�)B6q�Uq�4�j��YP`�>����L��:�%�&IDZy�#��ЀJ `0e��].�t�d󩪵��lq��d�\�R���t��?Lx%Jg�҇aUV�c�HwO�I�6���%�*����	��e�?Zo�e(������7l�y*��ܻu�h�;X`Ɓ��(�(���[�_�W�Ii�VY�J�&��%�j���S`g��C��G1�R��V��fZ�i�X>\�w�f8����-���n�t���{V�?�Ox2� g���Wuӹ���&��nV�8�w�˪8�ڌ�a~dfPJ���s��ġ��e���囜{v��KɬWV�Y�G�4��s�����x�8Oѳ�0���"����D����AL1�,d1��`/?5[E�y�."�j`F��/�ᕒΟ�9�����g[��:�,Ou�'�q���?e+�?�Rm�Ж�#��b��V�����z���7m��X��S[�,Rq��n��X�^�AVV֬���x��V��)m3��`cߗHb�R!z�#�JF��㨗PY�x�����	g�dU�lL*��r%�p��Vgs���A���5@;2g��q���T�G(2��#-�>� ��4W�vdlE=��R	�Ʈ�O���QPR(��
'=z�M�M~�Ɩ��ǁ���m=\�b�q=�Z؏W�s�ӷe�y�d����D�-���d�V-�NDK��x�,s�eu�y/��r������u	~vc��Ko>�8�b��TVk��w�<�J��M��H��W�L��b1�U��p\vM"2/��U�q2�R�]��Ep3ĜF�8��%|E�`�Ɋ�`�m �&�����?#l��͵��Nf���11�q�1.�9tyh��@�]{�*��[+F@"�*�^��a��x�!��8��(������wn��3ܑ��U�fS�O�	����[�,q���fM�R�5��5A"�����|����<�u� �+��P�;0�	.*���+����}m� c�v&^	Ep��E|��o�����9�Tf(k<��J��h�壔�J7���4��L'��������O�4��T����X��M���^�M/�Y�%|��F��PL1!wd�� t�3�TJIl��(?a����LK"�sy�?d'&5��`��B��_|�W!I"���	�.� }�����Y���t��,Ž�������H{�t}r4���*��� �F������y?%�/_��%z�B6���h����m���R�����f�Mnd<5�^\7��G���a�O��x�E[�m���	�	a����v��Z�]ru9�:؎����X�/�w<"-����G%<O�o��a�?�*9\2-mf<�H<P��'��X�#�L�SE_hE��3,�}@�k�H�v��V����J�C����i$�3����&8,��ƅU�)�/��v����fY�G�LE��Qf�_)�4X��W[�D��h*'�E���q�SyT��ʐ�\ u�W�`�8����Z��X�D�2�l�fƶL5��B|�y����j���I�&����*���%#/����,���7�c��2�Kܰ���>��I���x	�_�i��d��5GS�r�z��wl6~�6��r��S��D�z�n�=j�$�T�*�i�w��x�j���<W^.�	#wm/|��lTɘ�8�t��8���!u�_eGԋ��,��8ftqH��%пy�T�$�hl^�~m�gE2�"M��:�W������u���+/�,cGʝ3=���v8x;��7^�Z����/|娒*�����;͈j#�P�W��hx�G����Q�ʾ�[<D5���:�xf5:�X�Чwa��96�D�����&�[0Rx9<�6�*��><���\�"|�l$��_t�xbٚ��u?U��Iv�9��L�T�"�{v���a/������ߢ�������5�?�.L�[��PD�j\c�G䔃2��r�p-wX*1��Z�GV4㏗m�Xw�(b�1�O�e\��>Y��If�Ȋ{���G�lP^���,�V�ⳑ�3v3-�@���L�tF��ؼwJ�rov|�N��: �X�P|b��t�:��J�1s���sy+�KI�rE�3��p��Iv�J�XPK�㲀\���r�FjǶ���c���ۍ�zGN�>y���.qn:�cb����}8��t�b,����m��hq�Ǯ�C)��3� έ遇�E� ��P��5��*�E���۬�?/?v��r��q9���;��������%�7�TCG�����\�B��	�G\�P�ߤ��*��D�h</a,D�#�:�b'�Zi���}�7Nhw�6&W��u�z&3��/^�-I��Jz[��C��hW�$��~v>�)=�L�?29"A���`��\�Q�t���5�^�ᤣ�� 7R(XUeSm��s��!�����r�Mͯ8!�� �k��`�ͭ	��������V�9\l��^4�^�!='|@=�xO���I���;7g��(Q)�������K��;ę������L<�&_���pY���J+v���Rԅ�
�����[y�ydE��/y�[�|�*���~t�7�Y���j�IDC�{�}r;P���O�y	�Rr
�������!W|%��2n�ܫ�A
�Y~�aiq������m�Ĩh����m(u2�C�:���l�q�s���j� �ē���[�_	���L�l- A�eq�'��&7{n��Hf��;��'�;p�hD2�6{%ab�<�YQ���x�	���u]���zyx���}"�cJ*�<+Q �i�6�o�pa���zn���C�ڼh9�G��(N������`i�,�o�����
�k֩�K^�v-[�'���'{s���u\��-�z�VGt�U>O+�@d$�㯰�Zg!���5��y�	�U4Q����cdt|�cί|�E^U�d�����1�Z�x����~�26O%k� 2+N��ε���Ï��Bf=D�\_,�J�uG�}�TH� �ޔ�#G82y����@��`1amyO���8�ވ�~��r��_��!����3Os� �4�}���8���mZ"f��7�#y$�	ʗ��4l-�	z1�XIP��F\��fA8`�7}Ma�ܠ{��^]Q�ћ�&���a(MM�rMp�DY5�/}_�K7Y��c��2ze�pM�=�?݈�BR�3�ު�(�yy�=�"�����bͰO�0� �Y!�W��7"�2rE[�;���o�@/�y�FA��~{���w���C7	0n�M3�@�կ���w§z����;�2������\�{э��:?gaA�����d�p�����b�	����ڇ�qcHՎ�6��X��H~i��@���^E�_b)FZO-�I@�G�"�؊	Hf���w�`2�}���>xʫ,Gْ:�ox��ܹ�A�٩����ж�J��`&�hG�c�"����O�SqSx��b
@�����9D.G� | ��^��'B�G�4�[c��z'.�0��.;��k��+�ߋ>i�������bj��/��G1R_���H
ȊIZ�f��6�qZ>|��BC���/�{Hkp�Qn�>H��H�ֹ���׮�o�Ɯ�vG�>1�U ��j`�%�VE�������U�ר��G�z�64�ss9M[��y���sNd�^'�׵�ҙ�a�o���L��[��/���!j�Z}9+C4���z�* 1(�ڜxM^��|SFJogq
�"i(O)_5��2��u�4�]��n`����͉�|�2
w�W�y+
�'��{&��lh��U�D4�o�񕸚�{�������*w��`��~�O�_���<�8�/��Y;\���k;X�0vL��̈́g��w�"��-t9kS[}vx0Q�v��}����'O���,;��˴�>���w�d�܉3�x����/���k(��ӷ�3�A���J3�*P:����&���QHK�������n[EµY~�4�� Oa��Ug}�/���+zM�+�4
�����|��ۅ25U���zЪ�A6h�0'�j^��#YP�ٛc�nwA����C)֎�Q���e��^������8Ҿ���ۢI�v�h���y;�Ӑ��Ɨu%�ӳF>$΁����Ǿ�'j�'��I��
�ы$�mp�,�"}Z��mA-K�ݧ0)��$��4I�J�:�$�LʏS���۠-C�iM�д(��J��� �.Ԫ��s��m�Ȣ��9����FķA~NC�`��:?�	s��ڂ��0����,���K�c�����;S31���&FJ��#�F��E������mF�uW�y�1�P���ѩ4yK��j]
�ӏ�Z�_�,�/��.����͍�����1���b�2��-1��gt�����
�j|�ןT8Kb�k�XYg.�B܀u��?��hd��-H&�V��NV=ik��2�x�%�YD��x����F�_1���r����Ffӣ*؋��H}��H���}@n�O1o�E�{�E>Ѧų�D���
�E��4�!}x�F��gA ��4$p�*��.����2r���a&V���4���s��4�Y�^���#����hB_��Co &�unI]Qނ��>��;u���b�^?%`
-f��i6�s���>\���y����r�1Rb��4ԯ�\�&�QG�慊UZ$1̎`��b�μ��XJ��	����X~K֬���M�anw�"'�D�搳�C� "�ILEhR� VcVV��F"|�2jt�%�Q� �ѯDG����PQ��Y?�4�gS�L�դ�m�%�e��/P��	�*�zI5w�a���^DlX �T��RQ�huƈ�ZOu���2��2���V���
�!�}O\�Nj��/�_���h{���ե<,����Cx ����M ��J\����]K׾�$�-0F�B���d=���8������B�6_l9���ŝ&��rl�� �~���6����������N�p Ix�+@_�>���QN��]�+2�gxgeё�P6��W�=���"�o��Ĝx�q3��0XM�L��`s.����"?4������^���t:L*m ��l� �"�ɍ��w}t��,��N;���BЯ�P��r7mO�B�Ds*yA?F����º#yOg ��R�f�&��� Kb[ ޹x�#U;4�B�s'�NS���MK�;z�[פ\ces���*A��/�.%��w٭�������v6e�bǔz�όp�������Z�E+[Ŏ�/K(���4$$E����6;;g���'�𽏟�� �a�W6t\\�����v�s�*8�rبy�hg��!;�4�~�9�sH,��P`"@}�����P��yz�{R(E�l�����{�{��|zXX���#r��*��P�i!3�G8{�z��U��R���!��a9l7ǋ�������K����|��a�������:W�I00���A�І-K�jfaY��HB���Nl�~뀀���v$h��6f(r��;������iP�����L"tݿ.�i�w�R�3o�V�W�I��qR	�p��H���(l3<��t�f�6�
ܦXNל�t��
)Jƽ�D��:��e3Vf�����hN�����՜c�m�~�R|���;��1��"݅szT�{ۖ<�W|v��Z�&��c��6�S4���Pl��2�B��G�4�z�����G��EK��R�P�Eb��r��@;ښ뇍ɡ ��`փ�E�<p�|M���	`���L�� ԅn���8W1<#�,��;�$����O��N,�F2��������u��*���jɕxMDd��ٟ޲���N&o�Y����� t]*ϜM�X�N���ɒ��̷W��,FJJca��d�UCj�Q�T��[�ɮN�F��AhސT=�ܫC{:��Ap4�U"�y�yu�^RK��91��NK�6]�G�q�V���O��8x'nj�HɈı]�G-��'Ԍ�2��[�[5��}p�#��R90�u�h���#�nv���:��ޛ����(>��n�=1�7�S<�{B���*�CF���HD��)i�ic�nW�?:]��¿衿K%Ǧ�1o,�a͒�G���(�,X�P�Md\g�Hk��B��.�Ht�ĸ
'9:�������A������6�D�7h��j6q����>f�ku����1	jr+�tCzF��?�ڵ�%��3�%P��nC*F��:�6�w��/�p?"�I�c~@.)o _�2Z7��X�9��Q|��֥H�Sm1"+0[�)Ieܝo�
,[��dOd����|c?:g;=�1�&'�9�s�4�{ �����[P$J~M��Rx9.��mJ���h}L���1G� �����L]c<b.�X�&;C�7,Z�/�
�dQ&�������z��`�%Z �$�����a���T�'���QM=K�L����l�Vi�B�6
�a�'�N�lkۻZ��5E���^������	Y��6��e4�����R*� ��C�&���K�U��2���ge`�_T��ڗ�_�&�(���x�r������w��V�O����=��W1$*%X1��?�M�h��&���&>��!{�/6E?N^�9� =��p�c{L1aZ�x���f�+�Y�"`�!���a�?����I������^y���-n��ΪM
���sV�Hi�p��#��-{��e�I��-�����oA#��/,e��8R~z5�V����A<�T�L���
��W\��:+? B�f�d��d.���zzR�q_�p�l��Ν�vX���՗A��ߌ�h�ʌq��B�Ε����Z�E9���d�C��dG>����vȞ��9�c�q�w�����T�2��
�G�]u3Bڳ��Aɼ@�pu'_��A�Di~,�pw w�&S�ء X��_�Po��u	j~���8ho)���rhS���f�؈�� �7���^J��N(�t�;;���%<�
&�3Ā���&�"�5����G5��TGbT_�$�U��,�6�aإ���+��Bг���2�Ȏ�A�h��2%t���{����s����v���Ӡ����\ѝ�\s�K�N��_�����l��a�L�jDfl��O)k:�H�v�H�p�����4R����RE��I����9me���V_�;���\�o!N���W5��ccX"��U���m �H;yn( �$���]���0Ҏ�6�"���C�)�gb�$.�!vU� ����Ju>fi�����.���i~�7��V��}�RǾTX
�c
P'A�,+�X��En���R��2 �v���z;b����9{��V>�����mA�8QRO���[�o����p��4��ξ%W���5�<�r����Ӳ3��A�s��Z��]�}��z;�nmW���/�籅o��\���Y���PVl� �f�[�gDP�t�����]N!��ϔ��V�v�<�o�g~M	��O��n����پ9�I��~]袇�����ֶ^�T�a���2�����p�}�J39�����?-D #To�/[�P��\����+��d	.Vc��
[�h��1����"�4�#��)X�j�%s4�6Al�����T���g7���gN�����s^�����MU|����s��$�Z���Ж��JCo�7���ݛ$
�]�4緬	֦��<Z�r�S�
Q���L%@5Sz��S�U|�K�F���$GR$�̶���o����1m_ -ci-S�mr�0d:vKh�S{�&E"��=g�w�?x��.�֋���/'קG(J�(�X�C�K��Wd��ܻ��� �� ���F���\�B�t�c���*��Y�g�H�h������7�=�Eo'H�;��(�����ڤe���.ǹ<��bmj:�ͪ`�7�m�S��#]NЪ]dq��fJ{��� �i@=���Mՙ��_�mr��(@,k���oOۜ�j5������X�(~�9��劜6���M�̪*��x�;z�羇����6�'So>�̯�ʘ�X�=6Y��^� �&$���.�iA�љ��C�nfr�;�cZ	h	.�P����F���|��2:J%*�"o$�ג.8{�\ߗg6�]�QD���Y-_���^���h#V��d�˔�����4h�CwJw*E��a�
K��-�j��[�e~��v7�i1 ko�]8��E@�˕�]P�0'U�QRy�|��f&�*��ɭ[�%w�����a���K����5�@�+�y�X��8��گ��<�v<6������jQ	+<~_�*���#�k��7TDRD�����2�	Z��/�G��� ����bo�������*�<�$��q[׵Ic%���k������(6�T�+�:Ӂ��{x�`6)�x��h�,n9J�2viO��9�J`A2�g�/��@�^Sh���ʏ��	nI��O�\�z@UE��u��b�֬�Ǖ�2�t��k��c���|�`����Bμ��ّ�HE泣�^0���3c�R����4��F�u>���7I��o�"w'� ��*~�(@�_H�_&+.8�x��ԟء������49�e�-p�Y����3�����M
G'�I�H�Hﺈ*������Ř2�l]��h�J�07��͡�"�5��,��!�����Z��[�;�;gg��*�IO|���+TUώ"�s���6A��8�s�Z?9�a){=�0�·>����w"y�4�E�z�Q��
�Wt��8A���� ��}$-R#d2�A��Ҝ=��l���lރ`B�����)�.��h�`x�)���M|�T�7��� 4��+�����ᡄ�Cl�#�bI�;V�U*�B3�8
���GIh� ��f�����A�廙J}���9R�(�F�T,+H�$�0���Q_���U¹V�� 
�4d�+{�H�71�'i�e�5Qr_�t���F	�贀6O]@�C��8��=�K��M�<�����4rG���j����&�j���7���n���[W��K�p��� �m��i��(�O�Xp�S�n��汜���:~�-�[lJ�����@��#�+�'I���<�L��JH�"P�[��zUH���P�
-���-�X�B�����+�ږ��+�:��e!����$w���U��x�NBy;�1y�.4[��SQ�߅gC?������뼿9����l�r����U�n���vo��t��5���.O�[�Y�E�*���L>WH�M��O��u��I[Yw ʼ�\I1Pr�<�x9�9cZ`{��GS�y���p4`>�V�F��[I�֬�e])T��a�T�7���T����`sB�T�?}]ﺝ8?bfj�J^��0$NB7�?	���	��Z:�eW��h���x�`2����h:�F����x���J��>��-�į%]\>���iS*:���� �kl}����_�;�˧P�*�(,���?���O�V�S8o&0+��T��]I%v�4�P"���p�	��3�P�w4�t�1��ʵR���*�C,�=�<��'|2�(vz��L��3Y�p��1��	[�����ԃk�0D#� ��V7@[����Uy�I�g�6�/?9�R�)e���Ü���yw�w��)�gb�pe ����p�U�[��ol0i����+�ן=B2\j�n�:1
��5����,��)׭��S�[%i�>����o2v�o�6]G�=�ld��4r����>N;߼�1��n��7�La�s�#2��c�K�Gt���2h*B����{å@D4�2"6F@�6�~�d��|D�猕I�[y�Z�Ҭ}����P@o΢�w50�enip>]���d�Fbm���y��k��si;��ُ�D��c�����IY���G��Y�C�},�M�
I�faNP�:�l�{�L81i_@1�}rbĜCDaD1�����{EnO�iW7�ή�.�k
�\��2����Y�Yd�J�E����"�G0-���	��U�w���K�ʱ����NS;!�1��]��I�.����I�0�z�l;�:�S�"���	(3Uκ�Aˎ�/��⺤7�8�3�8��bA��Ͻ�"�M,4���+G��I�gGx^���!�:�B��4Ƅ����2�+\IlŒ^�yA�>*�!hE/*�fA�F[�Bl��q���`V������Z�<������VSTn$����Bb?i�.4ҩ䠪�O��D��D�ݿ�и�Ѵ�OӪ�10��	8�uh�Y/��"0�/,��Z+�}Z�s��Ze#M(��ӹ�Yվk�A��:v�F�[-?�p�j¥�,s��W�k��")۾��~O�������  �ȝ�?:Q3�7/Y^}ܬ��}lW�hOL���6���K��Ǳ�^���3M�����T�6��)p�gF\��&�� �#I�`������M�噞c�o!��>�Gv�'�*�����zפOu-m�yc��3����4�[���/���/XK�D�y��q'~���c� ��[8��Z/��I��N�u���n����q��+Z�k7���,qU���a��S��{��'I�5��@��{��Qgǒ�J����6�
xf���V�"�r��Ǘ�lؗ�Z. ��߀7m�O�ށsM�� ��m�]��-W�=�̩t�Ҝt��EmE��C��I�ZѮ3���0OF�y�Gw��t�:<rC@�.�E�-M+?��#|?�$qD��"J�=�q�*��6"���lt�p�_j���&��4�)�*b�b�=����<������~�/�t���0�u��W�y�X5-`i0,��,���q������w������D�'ЫBR-�\�h�	��I��`lv	�Ζ�X�;�h1?���2fKm�QP���9���w���s�ϰ�K�6���nU��IrE+�F�jG���\��9(o�������d��F0JG�vI���,@�����`���m���[F�01�XK�q��Z���Z�R��~� '�a�ps���V��7f�҂�V�4���5}��DkC���"��>kz�.����0��̐C!DM�,	)h���¶�G�h�P](<|T˭�&@�$f=�R6�d/�<�����~�����@� ̾5��"����L t�;�4'+��R��.;;��~j�m�DJaii��O�������|'�ow �C@,��nkzL���u*BLW�jCQ��N�li:�6!QQWe�|��A|�p��nIJ}}s������H�&V�9Y��<�5��_\Hw �B^�����񋋪֚�@m[#�����ν�$�%�?��f`1��s2\g��:�j��A߷_�9��b@�<s0+p5q��.�m�Og���IzՆ��fN;'��A��Cg�T��*�!��а Qna:���G��Hy�NsW��y��n�eRJ}���o��\���:���������=>I�Mv������o��]�-A�1�+��Z�u�\-�\��bW<&;����O�8 f*u�O�:
�B�實B��H���L��g��VL[��]�ԇ��4��_�b[<��q�j��P�`ȇ�=~XQB�5�"����/�g�<*r�Y��E�#���L݃Z�BPR�☢��g���ǯ���$��<�/�����т��i��2,�T��q�Q� �V���Zyc�%�8���Ӳ����\AO۔
 k8\s�9��mFov���ޒ�-�O�O�S��6�~p>�t�,��]m^��ۉ�s��HY!.���d-�,�l��|+f��h��������8+��ˁ�F��T�Zaէ��|�&���eAe�uxJ=��n�2B�E�X��1�{-��_���]��d�z�T����6wm�����E��Q�\���~L�d=U���Pj���y}�����1��GÂUI���vd[�ʶyÐ����d�y�h�b�?�V��e���4�I�.��D`}���*�$崏T(z1�P�?IpK�Ka�`��\Y=��h]/J�zr�(��#�qI���M�ׅ�X���Oo�h���+�ڒU�iC!��u�
�r�.I�t$���m��V��M�bD o!M]�骺�Zć>�rQW�&��8��9:�4k���\X������(����ʔvu��a���ꆋ�R��Zbߦf'q����a��B*���^8�>�&��n��5��H~���<��P�+���>}�+����V߳��pw?�v���I=Z �.���Y~K��6�j`ѥ]�<'ۮ�H.�:t
a�g�Zw茣{o�E�������s0�$�]z?e�<AjD�nq�qp��'����:�:&��= �4G�J��Q����H��c�6����Â����*N�6���I0�V=D��˴� /=,Lk_·�:Z�_a^xi*�uk�Nx]T�Qq��6sL�]Dݾ�U�������;>�
)�m��E���¾��	��\Go��~�L�nfU:��X�f�:Ob����)`�t�����<�HӁJ>fB�"�٤�'�]��'5	n��Q��O8���	��4�9�^=�;8�T�}���f>��s.�X��J���D����tIBӞ��nL�gG.�Ob�_Hp�i��;�mć
��V�Y �4h��J,���Z����u"��>�#W��{-�WEH#=�0/�65Y�s8�Hb�I(�ŇHl/gc�t��]�UP�b�4Q��3n%$:��������<r$�0(p+^i���}>��'`+�vo*#;�)���֑����q���>��A+�y���n!կ�n���vd�C�^W���^>��s����N����Wa-�������Blbю�7C�3c��>�g[I���^���I�-K5�|�4��0�3C��<��m	�Ж�s`�+�D�m�u|(?sψ��.ftrm�_ݰ�)���ͯ��]�y���c~@.�obA�Z�Ȑ���_!^`Y�gk����kK��,-��$j��"p�nU�.fΆ
���+#��v�?^|I���btq.�Kf/C�ty:�,��~��^�x6� A��mt<�����~�o�lrߟP�M5�gJJ�˨}z/`�P�kA��Z�(���;��o�w����^���r���?�cU��Bw	�-�!�&t����P��U�Vw���E�$i�Т�Ui�*�y=>7i�Z
���[J���dG�j���c�t�|��#v�5^��<W甆�ޖ@��ꀘ1�sg�3���sӲLVib$|�g�9�&i���>�<�K	��dG���{�.���`�g��XI^���S�wE,�C�������5XC;�Ņ���	{�;u�'���qh1Q;]`�즙�F�k�gҞ[��W�qZ���3�%-?OϽ�7�� �
ɍ FP꭬�2o�e�8��v ��"h� H�@��I�b��d�n����Tw/�+]�w���w�q1�����k ?�]<�~d��$������Z�0�^��'�|Kk�b9A��[%�%�p��޶�_��wQ��Y�8�"�Bܳ־t����z���IQ�јN�x/���zafp��6�t}X�)LE��T7d/�e����y����� �s���$��k�}\��Q.�p�l��e�<n��~�rj���۟�I��l�O� �4 �D�6�n�@��*(��*>Z=����q���"�kx�'��bz������ͳ-촅��&�sġg��]�'�_��H7gf�MV�l�a!�<<h�[�(�y��D&g�Q4�[
��;;�FOК��:��"`�KJ��vg�������O{�1	n��$3�'�5�����>%�I����ϝ���"��������{I�hc,|��=>��J?�����F��pxv�{D;��E{4ВQ=�c ��U�GVe*��B��.���Iļ}� f%n.I!;>xK:o���0n�@H�������v�˗�k6	<�u��ٔ�*]�v���1�����Mh2��dl$.#  e�G
�����jTqC����)N�5��*���H�y��*���S���}��y���+g�Aø76�o���~����dy݃[Ƙ����B��j���]N��7�3�!�2���@��x	��#��Y�μ���G�r�0y���~�k/�?� ��'�X̉��8}�8���W�P��WE��d�)\���li�~��S4�#B�nIm$�e�$�/�6?�����$eF��G����~а�V�G�S�S�׉kE��J�ݙ�D��@z�a���b�Q☵��*`���׍��4��-/^�T�\��I�O�����8���>*Ίo��dT>H��l��S3���1r��wQ����'���/��SE f��yWhU���Vc)˄��|9���~̖3���ټ:�4��G�Z�JC���ܾ��p�}�6Ɔ���1�B��q�e Y��\ޫ�l����a��w��١ĸ��.�w��kR�V�[���"�Y���A|�ص�^b,�VT��E*,�`TZ��$~�C����I������Ꮫ��B:�^9��OMu�Wl	#�[�*�G"��g\
�vY��M�nj�~cb)]�X97GHOK�TJ��t�P2�Wq�2���w#�I���=���E�t�F��q ��ϱP(�ZB���}�^�/45{�$,U� fu�w�Յb�<j��V�(s18t5���>|W��Z~�єd�G���%π�mo�d)?Rh�r�/f�5�E��v�k���ra�Q^�#c�7qu�3Ig���ӈo��8�f��9 ߶�z��}$�B��s)�|w�̿��eŊ5We=#g��P����7ry�7DYU���h�XJs�Y!�����߳f�:f]֫댒`��<T���+���q,"T�k�U���3Ŵ1:�@�l��!�{\��u�Z)uU��S]�F1�*W���#�Zd% �Y����*� +Ѣu��ȤR2"��1���u��<��˯�ـ�A�$�ܔ#A�1��;���nf��@�
��FG	�PR=U[M��?�WOvX���z�hO�~�`�w1��I��f]�|)0�;�2��uٍX�
��1X��7��ٙ��)q�3*zr{j�<(�R򮇮�+�>��sG|��Xz
�*��Mݟ�	��@��9x�$��7_X��7/�9��}�|:$e/�&��9p�26�gl���ޗ��$Z���>'#�t�� ��|K؅�QUb�}YeY��Ha���Y��ʜ���)U��?���3M[ʺ�O�?)�p�l�;Mʛ�	��#��bIVZ�O5����ڎ��E�Vc���1��q�WA)��+��8��LAS�A��
b��B���>}t����6�a���^H�����O�H��{�爒v�dHq"��̑�/�86��Nq��޺��[�o]�r����<�o�� ����\��k[����v7��Pa)���0�ODؠ��9�����/�����u�������0A�בO���8s�GA˖0��E��3����ƇKk3��DE�l��$E� �����f��#�E��L�$[8PTj��*�RW�8�������}��@����^��w��3�/��` w�N�=v|�Y�ﴕ$�yu<&��r)�Aw'��o�C�8R[\­*"����sE쾫#�s��@��������Y?ѐ��Ap���;�s�B�_���I��͊'�D��r�( �˜?�hY�0�ǩ����@��K]�6?��`�R]O}oc��k�.��� �����g�HU�T��Ӟ������}dVh���3C	H���7r�?c����)d�:p��;�[���Iq��ځ�[�Q��h3�Ʃ��p=>�OvG�-!��(��@GL:*+~�-S���5t#'ye�$���02����ʺ��45�;�L��P�K���{�N�	M��j+%�gImU�Xjw�͖���X�{�NL-�5�Lx��(�O����>e�Z�|��0W���i��w���R���l�V"�f�F��h��&W%�����r�c�R1<w]���'����B֕��z`�v�${�1�%�{��C}�Ķ�ZVI`��j6s--tx"��\ȴO�߭��p��-�2�\�E�`k�Ɏ��iG,28�k۝�b�G([_ʕN�j�8Wv���pa>✩P
��"�V�LY�Ro��p�_B�-�
��^X�47-���YD�����,ӕ.�+�vG+c����$�SƻY�\)'ZJE��ɞ��6L~ĪU��ը�hEߋ*��+���.aO�Bi�)�Լ��w5^M�"�I�]N��
MjЀ��_G�wR������}U��&��I*��>�$�����2�x�hx ctOΫ)=�z'���J,i�� ��G�E|�}�m<. L����hE���R��ø�v1B���΍*xɰy�nFȿ����tn�a�b	�BL�m뉷���Ի ?%����#E*�*�9-�����͇%�9��A���׷�%�_�fN�"{��8�ĺ�w m��$o
z�1���o����(I�Շ"�ub�~��2�6Z4�F|��cw�Ѩ�Q'����D���lW ic{�jsNoI��M����ߴ*%�ö�0m^O������ԛ/�a���t:�x�+3�`�j��Ɖf�^�	��xGδ�|S\�ں��J���sET��x�I9�Ǯ ��G>~�Q�gb��_!��Ǯ.��0�U���r�i�����O�&s>�iv��yUuu�l��<�-�6�0�<$��[k���A#�m�l�*��(��#�V�Uf��l�.�Al?��M�՞�J�Z�u٦fAP��;�.�ZF�T��j�����ή2��.þF���GG���T(j\�v��M\q�Wh�E����!�w��K��6gN'�0���o�V|�C����.K�(��;Қ��򉀼=�b8�`�-$�ߩ���Vx�2����
^��̣��#�6�$�Y��kp�ǄsXLhI�!J/�RP0[� ����dg�PT\��?��O�B9j<��J\L;	��DyJf��ho������$�Ɔ�lf)�İرi��?��}Ä�cb�����Y�d�=��y����+�=��ϣݔ~p;Pr�6(��ݜ4�Y6�o��OKD�s�� ���y�6��;a$p�^��̕u����9?����n2��"��g6��*L��t1���<Ӊ��uLGb<���������Z`@X~Hk�)�bl 0��S�7�w�r7���ݐ�e۹�+� κ������y��f�t�:Ig�n9��T�E*(�'����BJ~�Չq����ni؝P:%�{�kƻ�ɧ� ��M	�+>�[c�oZ�,�NۙGQ#.�?�α�{��NC���A!��T�?��s�GI>@i��a��Z
�?Sg�Cl�ѧ�0�u5���t ����	[��P?�N�P�P��79����1k��l&��ԑ�(g4�7�E^�?⡍2��Z��#��[A �&��إE-Z9��-�����WӠ��ٺR��k<ȥ�zx�\�+�K������΂Za4 �ҳ$�m�����\r���'��׆�|�m:�[!���#3�����*[�|������9��t@#����,�t�4lM��_+&��?Mga,���a�Fn�~��H�g�4�Tgh���p�-��n��~�$$l}�Jx��G�asȷܾF�MYEN��Cl�#�-��S�s���)��{��v=��<{?��9��
���!���չo\�~Ya��s��|Z�2b��
 WV�?x-�<��}�]�Ϲ�}<�+�����5O:��<��E3	�s��n����#����@b�S!��m��/=�)@tӦ�;�A��u��ݴ�Iw���N;T��*�N���ŀ��SQ�g\�Ηm�Ւ2r�8.��e�ҭ2�Tw^��n��F%���EDl󐊤�6Ig~��Q2KJ#i��N���e���_�B��gyb��EAՅZ���}r(�Eh?�&��J�ϸAh���e�R�̣tq.���m�(���׫��$Q��)������~!G���r
<�'z W�|'�O�qg��r]�@m��;���mN����A����h�� ?<�b~���$��)h��ȶ����{Ђd;�Y��Ǘ�����%��%.᧪�{���|h�M��0�E��\ݴOf������|��K�	�����@=5�Ixk���f� �h�\��v�������˰#�m�G�sm��}�y�b�9��3�����UdA~��o�O�<���N���L=T[��ĉN����Z
���R}�iȁ��Rˣ�`WB�b���T-@�̐N�ż� ��S`��E�\<Ǻ��0�qF�� �߫p�<���=9����a�T�M�Ǿ�}��]7 �8�u�o�oJ�B���˂���E�r��@W_~��$%Q�� 6����~*�		�'l��`\rm �;ag���j˷T� ������G_�4(je>���R�����pT�@v�����㬡E9�~z�>������(�Y��,�Ï,c�����L��W/J���ΫV�H�}ݗ��ܳe��WC����ɑ�sT��=pB��-<��I?y��Cn�D�j��IBg���!v�?^1���Hˌ2b��)��M��DH�l"Zp@o�w6��^"��a�[G2�������H�+�K=�����2�����"g�W���j�*N�o_l*z�C���>�ܣ��5a=�'*�M��2�x3@)	tncĥs�.μż
&���3��,$R]�pt/�.4o�9o�t߫;d���y9?n��5�4��H������t�Xf��x�����K���dE|?of�7���YV
����rr�d�\��bt>#�W�s���*n/vi�{�`N�6^{L$�a����ǋצ�v�}�ח�q�Y��{�&g�_��-�ԷoV��	�8J����$�f����uy(���x8BR3�uX�k\���<ː׍����jόA�r�BĕdG��}�C�w��:N.?�XS���{EH�䖍b������h��א��@Iy̎x-�����F�5��������9.�y����C�D����b~�"�+���F��v��=�"r�L*D��B��.�wڊ7���&�6.�D�k��>Y�탱��&���Aw�����GB��C�ј�m���X}�ob��e36�.���雰�5ܿ_z������m��̺ɇ*�)��$�؈���ԩ[Tr�� ��[�&���<?X�H'��C{1�e��W��������@r����^8��M/E�PJY�����d�ϣ�.Ct	�=v}��-�'�q��b(��{�M�Wa�?�d1'�İ���7�JU%�>�1������1w$�e�q�oڏGg��ݾ�/�MS��UH��T.��bZڼ����Qf�+������p�ً����H��>���IVIw��~�H,��=9�(d��iP�+(���G94?OR�w0�/�����BB��+:Dn��A0���=���( p@�KXOī32eh�t��3��4���+�i� Rh# ��ԯjI��@���
��a��P���M�.�����[����|Q��I��gƯ&��}o� o���]KJdxc YO6~�U��ĺ"q�DZ����ٗ_����݄F�u��<�-��o����aG��O8���	.�II�+�I�	�B�jV�Š<~׉a9�d��F�6�bZ]s��w+�ō­������R*y�i��
�~o@4s��d� {P 
[�1��zl������4���T�@l�q��D|�b��B��ݶ�i�@3&j۷AS����ʗ}��L�-B#���aq wު�Pj�)�� �@�X��n�}�t)�E�ssUyN���f�l�\]��B]d+�j�1a`�7V�(�84�pŽ|��JĔ�Rm�8yL�S4�>|3+!~W@=����Vfl����~)x��薡�"!������o�{�_�x���W����A�D���/}0� U�B4?�:�ߞ}pqT�+j^���/-O������&�Vl�=>?^9�n�-��F�:\���Q_���S�(
W����=+�(�{�`��? l#���n�ֵs���ڭ�{��{E��!�5������~#�K<�^�_�o	�ͫ��ު3eG%�N�v�9�x�l����u����]N�_S�0;0�P?j��ϣk�Ɵ��s��ꨉ�L�Q��'��8wr&��'�5���w��:D�$�F����2af�*1CX�� (񽢝�����P=B�I���+��|=�k����q8h�í�3!e�eUm�������� ���0�j	Ccd��r7s�ktV ��]�oI�!�qO#��rs
'P���i?�q[�پ�$�ŧ�7��G����q$!\��
T�OMx��Ws���sZ�uuYɁ���Mr��(��6�Km	�J13��%(L�_�����M�؞a�A���K�_�S�H�DB_�<%�`W���c;�:��Z��>w6w}*�Ly����t��'�Z�.��Z���2T������^�O�[@]��*S�x(��l�M٭�V��Rl�� R=y�|���T�W��@(�ڞ���������L�LL�Q�*��H嬑��������{ћ>�D�Y����=K.���+nf'u~"�R:	��/\.�`ĉ6TXqH��ikO�Gl�E8;%P��t�2�؃w���ι�&�w8��G5Ϡ�l�g�n?�� � �Ȅ!ψM�����7-ǐõ�B��tj7��3l���{9��uC� �J[̀���hG��7v��nx�"ֺ�%z\�EE+"�(�[(��~e�2VԄ�v$���Q�fp�L��1��]L����ЇV )����u `��~�`��S۷�����0V����c����wT�Y�����ra���}��j��̾j���r!�0_�o*�{�H��㚢����(/�RҜ��-�����'9�tx��4�RcA����ޕ3�����Fa�w���v��?b�۴f0�&tH̭R!\{{*q�S�J��du6ar�;�wV1Ɲ�*�Gq��t����ζ���{'ԩKPii���?�:cK���4�7p7�\.�����k$����V�d2}�8�i�@��-k!۶��W�k����Vꐔ)D�����L�Tߪ�D��3����vJ��(��?Ls�bal?e��s���@{�m�
�;4�|w_���d� �>�T�@t����+�xk�A�<}H���T��E�e�̥o{h�Q�*Z�����FV�o��zj�׾>��ɋ~U��@�bvݰ2�e�n6�އ6|r'�����A�ke3Bz/�8X�P��so��kk����e���Ngsm,t���^��M��P�s�7B;ĿߛN�M���zt��<C^�??�'�R��"���-FB������
�gA\��Q�9:z�Q{�p鰀�M |�F�
��Q��#*�
�1����}�2~d���Wiv8�9!���cS;�@��4��{����l�
��*��I+-8_�BH��ϛ�<���mAiG�s�(U��%:M\_zC{b$VOq���nb��޷�+��P#n����i���9� c��e�p��9Bj�F�«@S�t-�E/>��i�9:3� ��^�u����������C+�%�}�P�L`�3�ȭ\��w����"�#������}|��~1'�Pj�8<$h�od���R�� @����N���V�h�[�$=�,.��4�4f����N�P���&.��tpÃ��?��!��9�on׸0�!�"}1ϔ�nD�d�-vXm�ưɚx�lZ`I��!����}��0�D7z"��C�6/Q�mQ^n��i��2�����5pi�Z1�7�[`���b��-&���6�<ej�i��t��/M��C2sJh#+�wgV��A��ْ����� $�|{�ߔ~��=��|�{�"O�Tc��ŀ��0=�4�_�]S5B�Շ�<sG��J2m�����O���v89��e�~���C�zÍӤ�V�7�ғ|���pO\h�������s�ĮQ�7!��j��9)��i�~S��-`�QL�0 �h�����R�`���xN3uT��(9��.�r�f�%/D*��#րH>���Ky������b�}W�Q�;}\�Z9��ε)�>ke�e'O����N����5�Oj+��|����ٹ7ּ���0V����+9��7At2o����5%� �յ��gD���Z�!����Q�D�& ��ѳ�fq����R_�k�M5 %�4Tpo��Wb7l�6����=,ךq�3��p��H���j��k}�7>�n�U�x%�w���-(���,�3���RO��,N��=�C<��ɭ����r�g�(�#�E�B�귶ڛ�����.��:���;��[Ó �8��E�T����ޞXi�z��c��g���(�,��j�2���)
�g��6A��x�8��?�M��WNj��zQH�7�1%�%Z!#0�b/�xa��q�����4�$����<k+1�A�X��s/� ±O�+�*t�z����2�X�Z�c���_���J���vK�Q�S� ��f���;{�4U��9>\�z}LTï�Hp��e�����:-�x��iz��j�]yـ��/�fD�Q�ǋ��FR9X��_�	?�&R���I9�U!<�����Q�'�?7�QPh�w�Cs�40���W���d��BM;��OvXs@��d�1�t0���c�ک1G�$ND9c�h�n��#*g�E;Ǔ3�s�b%H9�� �D�g�y���D�ֱ5��Z���'������p���o�ZS^����Ð$�ja6i��@}��NBr�w����{�U����Ěs�6]U�����ʎ�	��Qbƹ�ui���{}�jӇ3�g1p� ��Q�N��K��1pH"t�b�w�ؿ04�-�W����^.B2��@�l�<��T׽�t���dh�EIun~?���;�W�G~�I| ��}
R���Q��a�Q{+���Et�}"�Aߙ�,�M��i����!߿�F
���M�'U��	�����^9�E�u&���"y��T=)����P��:�������q��wt���րU�aH��֤��hOYI[�q�,X:R	P���M�B> �>��J�"PN��b"��LG��zh+V�sl�֭ ��y�W�@ԕǂ��mc�4��&�u����~eg��a�!e ��g�z	��R�+�Z�s���T�(�˫<��
�Ss/6:�8�F�����_�Ҟ���T?�O �h�r�\\��iD���)�aq�BkTTSVix��
5�� �=#�`�i����].��� xXITK�TZ4/�U���z�N��Ⱥ�w�-}1� ��)�Z6�j��#]SH r�� =�9��t��t?�%�\4�B����]
�6<��!�&f�U���s�c����	��S/r[��٤�`�����(�*}*��Fp /�a�4�l*]j�۱M���t�W: ���t#̒�	��lm�-3�P��@X�2��^��������c$�dl�-�Ż�~�w(����{lˑ�h�Ё7�-ej�>>��u�, }H��f�7N�}q�2��6��o��e^��3�lb_�_!E��t�7v6��r���9�G#������~&�hPW&�2�~�#m�=�������ܳ���V��Jك"��Vg��?O��g�g�Q��FO���Y�s��k��F��d|`�f��2���s�Ne�6�gM�J^�w�`-��D�X�|��5�e�`@��ɱQȕ?�m�����cWzN/�#�IH�3�lc�Y��6�I�����#����Q��6��~���ZTA
�`B�
��%�����aٻ�{}�����k��CA2�Χ���S�=��[2b?x<2 �0n�Ԭ8.�M?��q�8�[=�����4"Y.��V2#���;F��䑾�澊f�O�Z��pD �|QaC��^��=x� �;�t���0�7����{�#��(~�9�6�XŊ�rٺ��)��[8�A%ye���Q���q�f��$���D��ls���`a�O�-'���>b@�cc>�*rX�Mn�8߭��ᝌ\��ň��*�K��wv�������N�S�P���ZS�.T��q�-�'t-��������?����^ɸ��հ܏���,��ֻavz=�מ/�$�	8�T�V�d�J��'8?":$m���d��z�)�'my�Jq�j ����6J�u�#ʦ�<&L�����
�f����� �T�E=��Z�l�1ujg&��w��G����Tf�6<���o�ˠvD�`o^�L �Rګ:Y�dGL�"��K�<C
�>�G=�o:s�
�4��2'�*�����<r6J��[���y5 \.�S*�f,d���W��h�~s-P'p�h;�7�֨�P�7� ����''�t��
t�ֳp�7Y���z�j�mq�1VާUY�^D"J�	��
̪�� �C��R����Z�e���M:�!��0���	"ȳPV�Z}�=ڿl�T�lBD���BN2P�\	C�(ș\�{ �n��-�����ݙ�ߝi�Rp[�װ$�:���P�o3�[œ���Ma֓l'������k-���Ν6y�[�K���FրqD�������N�,��w>��](8��I��0�`�3�ko�R!*僭7 �Az
�V6������:EF�`�p�����{5~x� e������Y�[�0�S��zQ���*T��8���$-�]/̭O���Dy�;�9�(��֝�P��n�{s��M-���d�f��K��?���j�����l�v�k���tLD6�8�;
���}+-�i!9:�MQB��̉����5�!k=�.7e�4ieܓy�JG��\�g�N�����j�<B-��v�����q��'�x
ڋ�a�"� ��:������ؽpi�Ɖ�*5�ǿZ~a�]&
�l�h�\��<Qa�3���� YB��/�bx�UD�O1��l�3��#4��"{l��^�i(��2^��I��J/�(������]�D=��&$%�K9��.���BSmѳ}HT-2jnr3Iz�yNY)��-�I�"���s�" ��܁Gp��Q��V�K!�i��)�N�*>����Vͱ�7��[}'"��!�T��$4*z��y���ՙ�Zg�vn
���[��~�a�Q�aD�F`P�v���1�UM���v+\d��G�(M0�Sl�6R�M�-�WJ�{���5��=W�N�֊��괕����@���w��J�dv�B𛪸��y���H�n���M�`�YZb��1 ^5�����ג]��am�#��I�h,:A# � uL�0�:��梳�J�cWa��r��("��[���߾9L�*a�����O��}��|XH��1�B���*���P<4����W'EvD�.߅��0:��l��ٹ?Gf���V�26���M�����[�$�UB��2� "fG��}I��yA��a�#5��+_p~^k�oª	XE�1�]d��-�Y��M�ӥY5� Q��4
8�q��Ï��9^	,i��9C��`�Y�8������n m0+�%�/MIU��7�>[�B���i���,���I V�_�l�\�O겉�y|~������S�߂ߪ{0�!߼
��*����'��3�>.��?j����v������]�ަ�ҥ-��=�e����+̊a�����L���0&����Ts	�S���ԉBA1#�M�Z8	�a����ꓞ�td8`ҖPk�VS:��hc�p<����f��6��N��1��MPncڱ�"��Q���q*���MFT@)��؜A�h�C�-g�(��t"!|p^r�/#��[s�j\��VRq��c�0��O߾u�#
����E��^�73�b'"�z�Y��#��*+g�� >R�>"�����+z������ZW��EX �J�]J���\���$&B���%��F#��BI�tZ-	����iF�5� �$�Y�e"l���(R]2�e�7ԫh�-��ڑ�S{�)}��f7xn�W yP���+y�꬝a�b�����3�S>�{[�Z@�L���'l�@9 ݱpVjb�o���n��@"��*��=�η� F�^�W�7�$�l�R6�:��|���_R����&d��a�ȩ�#$ZP�b�8dE��kf�a�I��a�k��Qw�N8͑H�v0�0$�3���gw�XD�M�'^��i`�,��j	O�bĔ��Š����g7K[X~[ӣ�a�m<6��oN����{34g��"����4k���v!e��
��ȸ7?����s�����ㅧ������>�f8�ӘY�c�<��>�K׾9A��Z��M";�	��`�阢��<&���{p���ҧ�/O#j҉�ɺ����w�R��5����; �\����b5��v�O�Vx�� �M�qI�n���!7��v�4��	��rv�_�cx�	�R��<4uM?�A5*R?X�	�V^����>��*�����E��&�1 4��1���'R�8�o��aD�2�2��}�T�HC��g��W�>�țB9���~y���,���7w��u6��vc�?��Jo�Y�0#���c~KB��H�s@SB�fǌn�(fv&)<Qi4��irci~��׈A�d�]G�(�������X��dSf�CA��yRT"�}��ݴٴ ��rl��wx?1�!=��4��5 �a79 ��4��[lg{����評��G3!=�V��\I�l[��=}.2�B�0^��>��*-�d�#��^��'��"է�Kx�hI����q�tR;������O����zU���|Ť�=��RŁ8�u�vK8[ڐp9��ō�<k"�/�kܮ&���$���$���LY��lW�����o��g͕�x6vߊ\����ɫT��r�1�v<%q�`�tG�Z"��TWN����.С���6/�#�c���hi��G¬�,��g�/I�-Dѳ���w����(7���$�DG���o��>N�ϗ�L���0N`��8�h�o��
�yZXo�o�t�;�3��йR\�:r���I�jH�.���i�^�\,�X	��1h��:���(Kw�N�� ���N1�bC-qg��쇘�F/h��˸�rv3%���w�D�f5��:�	m^Ğ��)���;��y���%/=&U �����N�=!ڵ�ݜ�n�w�5�]�7���;�{���y���vr�"x�B5X��e��R_�|E�Uݩ��!�6�IWV#u7G$ʵ8�&bp�6�9gsK�F�SC֒^��B�������?����5� �]��T���)Ū�W���x�{�l=�A����h]z��t=t4�Z�dĆ��\Ѽ[mMy�
 �-�>
i=ҩ�G	�Tv�ؔ,%�_�!z�|�R	��y��Ghw�@;l�P�^mh�s�4kw��C_J�h�p2���l?�C�Su(���Y�0߅*����8��6�W.���3s����іJ�-o�_&�����o�*�{ʠ�,��3z�0��6ՠ�΄N��i���+�� +>@�P>sk��g�8�����_����D܂��V,�հ":"��rU�,/��@�%D�%�����8�ji�O�����yUc����	r�w�E��3G�����o�9ōŻf�8���%Q����4Ԗ��#�'��)S��� ����� 	A��+�"�qP�����\��:<8frꄎ����K1�Yk-#sg��V�x�%�Vi�80�����uY���ޥ4����t�Q��/��ǻ��o��>'�����j��*+
�Q�w�<�j��W��Q<�'�p�+w�0�Kހ*�ada�j��^�H�z�8=��jF���\�A��&�&U�,��gkt�/k��R�(߁��&��4:&�G~�?����d�5APo}��{�Շ��X�WC3���k���4r�'�lT��)cq��l(c�l-��.G��3�w��@?��v[d�(�A��A�$��$�
��\.�f�C�Ҩ�U`�"��64�&}�8D ���[|d�C����	;�Rq�]j���pxX3��r��Ѱ�V��cI9���T�w<��@G��[��"�~����T���|є��El�9!�1��xK&�����X�I���ȯQJ�\�!;FH?������'��V���7��{��a�YCµ�P-{��Yag�ٔW� Ҿ�n;#ߌN�6c��H|�T㷮�k~ �u
�Bq��<>�Y��~;�2����<*�i� 
�a.���o	��>����"���1iz��;�{��^��~wl��ȴ�x��0Q�{������� )x�h��O� F�{�pfO6T����ރ�ȿX_�8G�dc��%� X�H��m.����<�L�t�τ"٥~g��D�	Esl2\ԲH�گ�Gd�9Y���R�N���u*Ql�D����o�������l{�3�����i[������Y8�[��+�N�OY��uC�|�5�C�+Ɣ߾��+�2����ƴ�\���1}`�d���U	���)���rVq��&ϜeX�ސ�� G��LĤSϸ"���~�<��� �uꈠX���|�f��=8��N�)���;~�E*�z�~�u�~ �YLG��P�eҳRYl���F��TX}�]���`�6<��d�lw�e�L���kT>���R��p)�#%J���vY��g�H�|R��	�y�}����/�p����2�3�w�U��68�˔f)J��.óKE�b.�"�TbJFxm�5{�9����_7�P9��s9/���͆M�_��PO";*F�	�����6�[G��44ob��j�����Ԅ�8�=":N��^�/}KR��DY�;V[0�Ͷe
zx�6��_�+��y�T��v���-���s0�#��y5����T���P	]V��XަB��*��V�>:G���>��І�H��X����X:�P��_y�@-�"����!O����qg�{Rڬt�'�Z�?�{�!�	�]�r��E�ض�����u�I9�����[�-���o^��Rh�}N	s8>- ���mq�����~�Իlg��P��WD�t���=�y(|���?�3[��4jC��ۿ;0�,�1̵trm�.�C��MuN+395�+7�j���5dG^�z�H�[Ëe'S�Ϻ�}���9��حx��U]H�β^������' �~��o蛉EA������m��O"�r'2 �!�^�%.�j�#��u�k��4��H�NOb���+ww�M��N>
�!��SS_��-�+)4�6�<�+�:E��6L�"Z����|GtA�i��4+�w!��P�[(����x��d�����Ө÷�2[=��������NW٣yc>��e
ӠH�aO9���F.�f��&N��{Dު ��������;Y�=V�B�b�x"b1E��@��q��j栰��ңm�l�ok����jܯ���Y5��Ve`:9�HSKS��-�?�dY���XE�P)�t?=�Coݬ|H;�JkЎ�_n��tz8ú�&�׶K�^��H�]��d�|x�g���,�x�=@�4m����M�=_�ʯ��^<5��+�xSLj��b����/U�8�>hT�RD�	���Jx����ÊL-P����b�"��Tv
Hhߦ���[A���`5y=^.�H���7ep"��v�U�0�x����vq75�x�;�T�-�E����_h�ZCH���q&�Fxe�@�X���w#/a_�4�E5'�AT��M-S!r�Ǟ3� q�����8����/8�����������̈́��]��a5*N_�׺�s`�~_)�����c��?}��$�c���Iz�[&�*�g*��	P-���Z7)�@�8L�P���*��0`@�KEա�W�s�HR��3�p�[;��:*b*S����r�-���g���\��$�/ z%cҗ���E]V��׍��ĸf�n3w�jJka�@l�k>Q!9jtҴȺ,ֱ�̕�̴��wPx����u�D����T��?C!g�J�^On�*X~��%0*�`����zq��u|�ۅɺѬ��#<�3�>� �eT�θl�
���s�$������9�Y��x;�')�����.2����Rs��6cx��Pcr �.$#{��6#G�?y[oFqu_oل��F;Ts���?��
�)O�0��4s�ɴ�6Cb�I��y�?]�t���e�Cׁ6�Νr7�i��}�Z��������I��o�jy5�,�аa�PN�$���P�ϝ�46�^�C�]��h�0��M�m���#ڛ��#�����u_�ߖE����0u�R_�iH�R����5V���X������Fћ,_���#'����?u�C��	���ǣl�W��C�Jx�^��y��� �=�����{S���f<��@�"/Wi����h!:l=��^���3!�[�l@gl1��L������K�\5�/̌�X�	�����O��>r��]�㪍38�g�/�r[;^��f}��o�����hզ��S�GnvJ��Aq��B,�WTBt��,C�_�.�lB�օ�%$��d�3)Ծ9[��Ģ���-- �T�wQ���F��lڌ�ь��ZP\�_���10�mn�1-�K��5J�H�l1Ôv���7U'��K�Z�T�&B[�E=q�gX�%W)��w�J8���]#���L�B��4��ǋM�ѧl3���@��#l��\����%/%�!3�`
ܷ�F�_��i#���}�{�/r�ct`u�D�y�3��8���}��U>�Z�\{�G�m�g�-̈��.5]p��w��:P	�������(�������s�l����pyY�W)�g�a��U�p+ 	�v)�MU���5��H9�e�`c��������E*�3Q(�-�v�}!��衭6�CV���4MgK�`��|�0�-�Y>�X	ܖ�$�����ɴ �k�w��SP���)��n2V�)Q�QC�N���e0��J��%wz������H>qZz�nv$I	)p��XY���an�ց��s�p�]�	%�G����xظ�?��7�pmf��>x�(qM�|�%϶�eq�����m- ��h�� C3��ȃ���,�ĸ�����V�a툙�T��@RW�|��%�^ ��
9Yn����@�in&[���1-��:V2���4�'����`|S3��e�߱z�����6�>��g��3������B ����S�"�I�>d]O�(�Q�����Ѿ ֱ� ���T[�l*�A|�$j���6�Ր�\J����$HO����ST�ʶJ�
2��hI	��y��Q������
�+p)<��Q�'i@�uEb�F`<8�q�U��/����w�4`��KD���i�;2E�*z��@6�aî�o6f��~m��M}#Y]�@��� �����D<�zu���@�̔-2�݈�aj��*�<�DJs�QדT�)i��C>$E��ɦ����ꮒ�.%e`�:?��V���o�PJr�^k]gǨ	Ӽ�	���K$<���X8��d⠶?��4_`;��PRq\xq���3�9�#@��(ŻK
	�?�j#�����Ff���l�߻363Q��u���z����1%�5�Om�`��O*U���^1ϙ������X뒧��eS��as�@�{�-]z׭�޿�ӣ�'��1F�M���t��� і�X`��0�әR��͋ƨ���!�7�^R�vX�&U�M�F���U}	�zrIv�Ka��(I��4sܹ㰼��{�Oare(W�wÙ�좪�o鋉�K���"fk��M��,/r�#�ݕݿ��ƅ�T<�[?���k;p,��"���t�N��taUb�*�ƙ�,Ԗ�x ���2z����ǟ����5��N��7Zi�o���iFj{2v�a��/��11�0jTS����:�>��A�r�?��B.�e#��E�G���E-�w[n�J��+%i�-}��?;S>���K��E�b�[� ��yb��9����YW��>VUq���};'�o���܆�^���)�Z�zu����A�v�B��E�%�<;�&).�`���_d�G8�s� �ڊ��'o�oqS`�H|�ש�Z
��j���P�9�:y�gwݲ�f��ka��g��F���[�<h��}�a���V.a���/1� ���-z�佌Q�UL5b���B{qA�e4(m��U��?@L��oY��'��2W�=+
ӰW'ɢ�䛻t��opB��Qso�o�D.�Ot���w��θ�6g�jZ�"u��%ze2;D� R�R���#Lg�?f0:G2l�x�+���.	.����l���-������(�o��u9j�)P)]���;T�6چyr�+l�`�gʼZ�sj�'ό��@)����Y(~�mn��Ft~&�(4�05ݦ�)�W[ܝ=&�G��OX/����_�.EBʫ�ς*ݼ�lim^t\��q�r���:�F�3�γ@_U�pFo�Я�9{u���y���Wy�⑷��/~�5�]�ҙ��\>��QW��g�"�K[���1C'L�!+�򇣽�lW����]���r�eY����ָ�-T��3�y�C�DK&,�O0d@D�-�5�W~w���>����+X�t��^��4]�!����zt�SZ-8��s���+����j$�"�C�d𾮀/��e��ol��5�Yq�ˈרF�3�m��K�{L����
�F1�%يW��A�� �Ce��҂+�rxݾ "��GSv���O�Ҽ &��׽}�3"���KƊ� ��M}�s�e}�v�o�Z�h�:�-�Z�2X��jz���������Xv�
SaSO��&һb�(h����ǉ�ĆO�*��-r��!��o�Cr�'��Lw�="R)�_��U(߲~	)�[}b����,�on��@4b����B��ܳ�W]R��_����x��/ĳH�E ���{����>�Z���DS
#��X���}�B\��>���=��rU���ڪ�p5���J	��EI:E1^&�FI����,�)���A�!K]�p����i�<
1tK B��D�)�8͋���tM�hG��Zl����.��H�=�ҏk�/|8�l�?���DA�.Pu��pؿ�bm���oM�˳�A율��Z=�߮�g2h��$�QƄ4�Cq�#h�GL��v�jfg�?�O�`�!c�!PbDj�?-�b�~��@�53^/E���|{�ҹ�T�Q�j�����'ċ� �5��>�䚨�GÅ��BGq).ղ��zf>���� ��~��n�!(�*39	�F��6�	���A�������D���cH#����~�b��Ւ��[|9cY�W��OMkZ�������<%�j���Z3��$X�Uu"�}aB2������K?��\�)�)����ȼ�k��橿u�]5h�	X�J�Y�X���2���҃��㬤��_��y�{��xGD�T2��-��H��p�ILR�e��ۼ�v�?���H����b�F���[l����1x�N1��r��$��a(*d�į:��_��9N��X�G�3���/��[w����F_��y����mս稤B!��`�N�}��[��%���Ԥv��Q���4�Fً�����h�����y?�@{,��&�Q6<�D�q���e�!q��3g��9���щ�~���PKm�Wa���u�j��j�,_�z���q�3�Ԉ>�@�']ُt��:e�I4�̦H��O�eq�a	�x�Ξܗ?�<^R���轇��_	���8�T���"�b2-i�>�Tr3��̳�;�e��"ؓ��x��,����\ɟ����-��z��?�J���=�l��>�|�����1G�4%V�9%�ME��&h�WM�jSl��E��5�����N�j����}�>��� ^s�D���
n���k>mÁ�D�Bd�X�'���>�R�v"�I���K�������d5�ݵ�nه�,���!����,�#�"���b�$����рҸg�t�]�%�����+4�����mU���u-�!CM��ҿ���˞j|RKf�Qt#�T��c2h�q^�C1!ex�,#.���f�@�Y� ��XϛnCE��w�۶4U��L�ˊc:�p7����_��ԠL�6ii��劻�tPG}JTxwu)7�X�ͽ�;��ys�cj^Q��-�gdڳ��l�w���$��U�jf5���ָV+�� ǒ~��|�M�W'�쿂����Lj�f�=��V���W)à�`�61��=q�g73@КZK^Zi��Z<;rZ��@�}�'�$������T1-T��^EQv���2�M�֩�U�D
@i\K�S,���R�PC�ګ���󤝝(�v�����w=��Z��(f�繣�;�'��֠�}�6#�*�	���L�JG{���P��zх;�⹫��p��n6Q� �&G��;L���Xc�&�Ҧqvɶ���������಴`>��v?�I�@R[�"K�ꁳS���L�)��` �*_�_�>#�g�CmJ7�bs�=8�Q%�����4�q�{�e.?�Qd�1M.���*�Ԡk΋Q��E>����_X�/���R��,�w��"Q%�Ɲ�؟������d�-{�ǲO�J��1j�'��@��R
�į��pN11t�m�h�'q�=!�#��m��Fir'U􅰣.��-���RG�k�_�j�k�>W����/ 7¼�<<�����(���{V}�Fൔ�_��A��%�-��$�s6YNy�w.�X���?s�WC�FY���!�����lGMВ��{�M�k������#��PBM�?�P�-��_x�cd��I��:j%(v&��k|*��L���B�\t��T�ӢsiP@R�=�D����[y*�ȫ��p����()}����.���5�w�SЃ�ܓo��1�-g�)vS��r�������.�&d�%����|���BG��ՓHd�1I/�/-�$�w2��� �&�1ǒr�b�#7��-�[�?�S�Y�n�2���V�ŮU���/�@�c �j�p�ZP=`�^hB��°(ĸ/1�s���lؑ���:�h�R,n0�Q�s%�趙�y%8��~o����:�A, ��C�X#��3�?R���%���3�V��#"�;2Aj6�U��z�r=^�P���dU��D�wcx�-�6�e�x�f\�nU߭}���b��ķ+�;�^!d��5	��8�h��A�Emg ���h���ݙ�x1���׈c� �ǹ3=�Қ��'� a�8Be/_�L"�/���!O�"	�՛���L��O�iO������͏#����'�7~��\|Х6ݙx�G���	��E�In@�ub�Z��jJ&�m�K�~U���OMO4Kcf�;��F�7����Яɗ�U:et} G�!�<�6�h�����HR]"�b���Q� �0�AC���u�U���y��%�
ɬH�r�s��d��8W�`�;��hv�f-�?P�������VAT�=)�+�4�t��穨�����Ig���#�c��e���O�$Պ HW� �Q�'PT��P�������3`�Ezf�sB�[�]䛔\����S�VJY%'���(5`��:X����I�'#��:^�Rי萬����U��n��w_a����r�-E��.��k��猋X�7���k! �a�����Nt�޶��$`�f��3���f<�,�#�4|�u>^bw�I(]l#�����?E�V�̠�iή�x�F�-N��u?��3��k�n���͞Ȫ�A���Md�(T>�р=�Dh��cً��%�O�v|e����x����VY��K�w?�B�\;;��ʽ��t�	���@��� {�b�aQ�2�a���I9,J2R�B��C�|�M�c��rJ��h����0�d�&��dGhOj�jn��(u�^A䂸����_R<:ho���0%G^G�\~S	�wtf��(Ѣڽa��p뛍~t
[?ͯNNC~��6!�si��s������~�����T�[p�;.}q�]�d�,�l��l��DG�9��JBJ�9j4����o��g�b��HK=���`U�0%�#�V�'_!X���AoA�g�T��"��I4#S�^�e[���"��%F�p����V1Yg��*�=j�Ʌ|T�.@���>~D4�ny1���Ϥ����OF)�n;~����Hq(I�,�L����^���=!b�;o\I���F��w�߄Yc-qQtB���g8c-$)��)�*��pE �*_�����۬�Da?��R�i�Y~�ZL���}�l�%b�.eH��eR��!(���*�$B��}��d����Tizڶ�'�F����$���oߕ�����I\�s��5�ď�[1Td��wLO��<��=�{��b�\.	��%�d?�A�N\0-ۏ7\�F|���*�~�3Rl�e�dl���hxU��]��jp���vj%ay|�&��}�q�_�U�B�N)��ګ�*"�bZ>)����������H�ϫ/$نQ�(|�G��+3�u ��������a@��b^�����U6)Mp]�f�m�	3����N�/n��i��ӸZ\�[���	�vA���`{bcRjC|ڟ
��q8nu��;���"7Q��.�Q�
���r�o�T��,�h��BWqW�+_����_���hC��ϟaE|�Q��F㽫��݋����,RШ_"�=o8dߍ�ǥ�~�R����A��3Q�]4�Т�S������AF,ͥN/��!ַ�$x�牾 >��*~�d(�L⮈�����_ d����]�zP(Ͳ���s���tش�6=@<�%'QK#-b�7�eHr2,�	��9#%��>j���0�^��3脙
�~��-�<������D<4����*��^��5�E����h��&�	�{���Zn.o�������bM�j)�Xٿ��gX�f��Ϛ	>=V"c:u�T(19��� �>C.�B9&�\��0���~1,K�|Pi��I��ݱ������P�	܋�r	͖��@�DzO_��X=�U��.����f{7w�ģo�'k3��k�Є���K~O���Zi�ơ�a�A��2>�����F��tp�Я��~q�298��]$�}��l����|���Y��T��6�+1�B_�t�W׫$�RR�� wP�0x�hB�	G~T
���0Q!�v���G��Hh ��)�q��%N�<�.xZY��P��FOU,vtT���/gKI:ѕ(-D�O8l��u�:;�J?�'�f�Uʽ���XK z��d��9P�v��V��(����Z��5��A����Cb}:�I(��;M �i�u��@OЙ��PK��!�Z2��)y�+t���O��ZZ8��먽�o�����l������@�j�*Q�#�}��"_�; ���l��*u��.�i��BL�6�
��Y�v�ˬ΁��	�}���vWy�X�Mf�o��DHd?�1�6$y��I- }�\���ϯ�F��`{�.d6�vt�_Wc��S��+���_N�`��
�m!�ޟ6A��>R`�q\ܼ���ֽ�)�=C�9����2�����l��O�f̿�Im�y,���S�#��n�p��E9>^F8p�� X4�W�m���p���1�U,l�k`��� �1�%~ENvV���h9�C.,q�|o=�h�+�p-� 7t��^����y %B��A��PIoz��\7Q3���i�K0%x�1���^�.�Km�/�3ƕn '��;�YA����Z�o+[��D��FQ������ i�<�]S���G�.�t7�H�6���rT��������0�������-R�q�.��8���]|B4�e�c�x�ڒK��?���G����7��o�~D����gh���:~�+��%��['6��M#7)��HT�Z՗7c��ͽ{R{�r΋\�Mh.q�@�-؇�����$��T�Ʊ^��eg�z�L�I3;�ݼ��:�"�!?��d_��eϩc%�����n-XN3v�z8�P3�������L��>�N��7�}O�!�n�+��\ljİ�ĳ;�}-��z�d��n����>���"uu:g��I=�ų>�+ �Nx����@�(#����42*p����E]�/'�Kx�����Z$��׵C�6M�� г�/����oB���K��/��-݂.����sϺ��ms]���N��Բ��?%5��b��ʦ�f��y�3��'�B�v�Τ�s�{A�|����~S\��=o� (�+¶�ߟ5����5�t��7���s;ڿh�,��k�C�+0�������F� K�����Ļc�<m:.���4¦5��P���aK<�S��o4�y���X��gc�9������>�����pǶhB����J�A�P>�#rd���(ED��s���O�Q�<aǕn�玮��r�w���0`����Ԉ����!+�R?M�j�"�c�<�j���GjQ�&�y���
�5c��B��L��6�K��i�*���[!]���Pͽ��a��S5����w����ԒŶ������C��A�W��W"�	���rާ��NÙj��;��~�G"���Y?]���a�~��
Q�)���|�5-%�c&�M��|@���ƀ�(�p��:t�W�z���� `���*|
_�t���r��w.%��9�g��$�r�	�سB��eH�>*4�}h��������
`�-�6n{c�Y�_�( �Y��9�'�����z��}¾ʗ��_R,��V�� .�� z���x~8�o��'�ne�y< w���*�h��T0�^�Z���{#����D"�6��Y�$w��{�w%�9bO&��p{f���d;����I�ث2"`�9h>��t*��3=?�"���u��mV1_�?�n����a_�
Mib�pj|_�]	Hf������B�����ZW���v�X������9���3�OI49�"5 &�q�'O��]���T�S��qv�.�&_��s'F��D7�]ϸҙ�Ft6��iu`�.�I�s��"�^Y}a[���JF�Hè�?<��4�]�@O�G���=x7�� �k�s��'�i{P�s	�|i�
�b�/ w��3SO�]��ND�ǜ�����Ƭ��{Ɓ����7%�>�y�Ă�f,�Kν��hLQ�:�K������%��A̱d*�bzߋ�/\_��}.�]�^֕�c�I �͐�e�*X���iC]B�o��?�� }]�8�w�Y<�l*%�f6ڀ�$�@�S�d�cd���Q���B����S��CKݢO���b��9�D�Q���9�
h�M�� ��Z:��2y�-#���p��1��_fiS/O�L &��"�����{���2�a� �5s�܇e�fژ�����)�@��se��u����p���[))��	��j�Z��)`�ɰ�i;E�Q��s��j)	�O����n�]������u��1�3r�Q��X���ʡ�VJ�n
��M���_s�@w�[3n�{��އ'���G\���h֌#���݁򊄯���yJ я�6&�n{Gվ�t����T�9�QnY/�p��;�_4A͏��F���g�����ǈ����#@�0�"��aS�%S4S�ӨBl�G⮆��P�/s�Q���;�^���ұ��`�@��
���>]t��5��o!X5�w$��z����?�W�+b*����ҦP�����T�	�6fC�d"�^�閔*3%y� �ꔞfo��#�QS�]�8��=(�ۍ�?��T�L؍yq'�AWP r/
�12'>��DΙkw�EW�&��c��:�1�D��ӎ��:�ѥ����OP>� �ܪ8�$��`R,�Q�W�OeY1X�����h�0��?G��<>�t�����+��~���i�qϳ"F���f�6��8`�Gt��h[>ض+���Č��Aݸ. ��&i^��ly~��]��ыYtpl�z����!S�S��}�V�"�?.w0C�s}%f��Ȥ�&���b[���2�mW4�m(e8Dm
* �$�ftY��c�lgSd�<���8-��3�&]e��^�47,�a���
��/t��f6_W[�� !��9����Ӯ�� B�\�l�n�)�dfT�q�uVx�U[�-���� ��/n��g�Y>������{ISBm8z`���N~�CB#����Z��>U|j���ߐ�fKKm��qb4�DE�˯�%����t���whF ;������2]���)�p��\�f&;���
ֲ�f�x�d�r�
n��>hI�=��]`�d.2�����Us�U�+��<N ��ʳ��Eu�B_ei`�.�"^�(�k��*C��8��$DKF��6�~�3�Z�$�bpiIU�?�K�[��-Wa/�/�A�k�L�b�G�#P	D���3�%����ġ���2���W0�J�oxU�� ��0<"��(���W��7T��[:���G����X�0d�{9ؖDĕ^��W1N�� 5��	i�q��T���=M�U��?�������4@1��l]�7x�)@ۋ��L�ސXGB�F��S��K��n��0��Y����"7�,�B�'���.���a��F����՘�ߨX�,�.���)�䤢��V�1���jT���-!.���垯��v7�����,�j �ekA�
�;Ɵ���o���$�� y?bѥc����L��e�Q�N��̔��=��V���RB̻S�|D�4~٣L�Cԑ^L��b�*�w���4�T<���'���Ϙp���������	���3�(5X�  P�2��� +c1h*X��ZU�������q�4މ�0R��>.b����<�������*rn����/o�HTu��Я#s3i�M�
�5���6��;��6��R������8X@Z�͓��N�U�U*L�Wy=�t���NI�@�L�3����>���ӄ۩�L�_�]Po
l �J�4Q��;:0�
�M���đJ����ؽhY��Yh�r�.y�Y��h��)a���2@��E6��Pڞ�
�nJ�wSfht��Y�c]�_?D�D���&���jФ�t9ٶ��:�>qx5|ﯽ��:R�:��)ƶ�ҽV����?/�G�AIOD�&���	�����H���"�d%�Q����혘0���JC�ȅ��&!���2�����R��B�@���p���!/r�7e1�����������%�t贪9����+���X��Mj[��E!�w�桰���@ �:�@>"Ĺ��h��mP"�n�uVt&����ș����'��7������[a�>o�r��1� D��c�C�ი��2�I:B��y)�&���ö�UZv[L���3�`i� ��ڲ����Wzu�L<g0��ŝodm��B�s���ӷqM�+yq|	�n}o*�����ʪޫ�� ёP�ji�!ƪS"�;�� {O�Ͼ�ݭ��9sѸr�l�a��
y�ع7O"�?���x�v-Q+L!<�N��r{�1�X���S���[ώs�e������	����zm���|���X���>����vSd�c�㣓d��g�OKX�uHZ��@�ԅ���e���o���}dA{��jS�_e8]f�Uk���2Du��g�>I-;�8I��ݸ�)C;��UM����M�5h4�V��W&��HW�a��~竵���sx��Qð>��̻K�S����\�V6f;����~,�����r��~k������C���F��DYe�w?��N ɭ����0��f���Sx�'pU#W����`�y������0	�$~�0׹��r4&���|;���ńXM��<�V1�ܷ۱wu
2��)�K+�k����&_;8f���0���2�2���q�L	�y����<>����?[��w�c�������ۛ���4��|O^~�,�
� �U~ob4}=`_7�+)J���_@�!��$B�fLv!��n��d����g��^S[O]t�����d�0��?�|��NJRJr%�	\H�%P�TT�f�˒}�<6�-�Ø�g2eg������%�x	{�:�U��, C���߉*P����Ua(z*Ś��Y�Pm��+�`D~�����k?�j�@r��+��K�J��7�qԹu��&_''�߽���Z:Qӂ���)��}���K�� d�t~��n���oe��FB�*�˃�&5�f�rI���_�Z�rUś�Ľ֋��]^k~����Y�E�(���{:w������֯zwE�#	ؚy\���Ö����Z��?Ѷ2 }*�Ezh�"H{!�(��4I�q�\p� ߧL�teܚ(�������e���:/�p v�mi��6e�:��l7w�'2F�ʤ�ag�{�<s��T&�j���0�\0S�Vl��Ls�s�1�k��b`T��_���Mk<�	*-w�
6��[<)H��h�c�V�X�i\b�)h?�3"�?��g�0���X���tc%4��L"`ģͣ�x�^�;"�`�#D㲎�y��`<�����W����.�7������hW
m�f��A����3U{�ZNB��Og���Ѕ�㦫�Bm�+����hs�\����0����+��vW.����q_�b��yx���Y68��bg4?�sS��o��Y+�s=Zy*�"O�@�B �9��Ϡ�^+L������t:�P�1q����M^��G�Ҹ<Gc��ÇM���"����9-��.-��E��Y�d�\��3s]��^�������ێ�Gf��`���k�VJ����5�hxR��6�o�~.�n'=�5q���m������/���ekj���HLs�	�	9�7Ω7���R���>�����]+�%M􏘹�����uoy{m�f��Xs|�SmOY�X]�ZnL�a�M{k^�͜���j�w���D��g	0
"�L�f����C�O��Y� h�!w���r�����eb�D�X&�~"g8=V��#�q"�K�0���MC��v`���<ZIc������;����ӗ� R�@�Z�x3]"n9������J��rk#��QEΙ 䥍���JI�����d���&�a�0�Zn����hӺ	�9|�2�(�K��AG#6�)����j���^eW�& 1.�gY	G���:Ńa�ʴ섷P��RE���O�~��a��r���	6,�i���x�t)�퍺A (�~3�.A��1V�I���W�V�ڼ���t�q�v�7M��ǽ��~�R�7@���Y���g4��| v1.�*�)K�Wm��(.�H�1�j}�/�
`�,v�}�r�W�S�"�اLZ��+S��W�A:�b]b/�����(*�0�P�T����1|
D�*��k��o����ߌS-�Ƀ(�*F�^H.�*���F��|$K�|-՝^R[1MˁFitS��K�S�=D�������eQk�[pd'�j�ⰾ��pw2U0ݞ)cn����̏���M�P�&`}Jz*�����ص r�^ߟM#�IUWVkԣ[��YR٪Z=��N��?�`1V��C�M��9*e���y蝧Y�_�5|�◗�y�)Ӭ�|~�r�Ċ��y���1�ݹ��b��]!5,J3��HEޠ*z���D�u��@a���Y38~Tqf��0w_~%7/V�yKI"tP�'����ԟ�.y<�y#�BZn��|��ZÛ�5��m$�s�!���o|��ٕ��ڝ�I�����'�7Z����8�Y��(����rSeZ5�C-?X��[p6�5��c�eS�u�S�$2�Ս�1�N+��6J2�ʤ�n�7ķ�VʓW4�������%��2���c�W���uqe����7��aQ���w���}�N��_/�J�Ѡ%,1���Y ���"G#�
~�n[�7 F�l
#0Zm�*f���y��l(㴷Z-�<`�h��f[>�N;.�/9
@�+��`',��Z����T�@4j���C�q��p\ǥ�"&���7��á�d��᡺�@e>t��6��P��S13�IM�z$G��V縣_>Ӓ��Л1˞)�rA˪L����,�7$��Z\�V!6Hl�.�Ez�����,+s�������IPV�^Y%2#;���c�%}.ὢ8��-�W�
1|X�<����8��@��O/�q�����Z��e��qC+��M�g(!�d阇a�����Hi$d��!5.��/�����T,��
=�E3 FU�'C�N�HT��,�l�Ay(��82�Lǹ�{�;�VX��&h�p�W�o�bF?v{V�2A�Q���a�Sr@K���w&M�M�ܱ`ũ���+�@�Az=�%�U�rg���, �2ό׷��0u���3����e���̿��(�0�S(ט�k����*`�]#���"F^��L�n24��ƥ�Tu7�L�n7,sXc��U����WL'�4�����n�H�_���u:uc����CT�?�DWa�bh�}�nE�mW�`��)N=|K��9�j'y�� �es.��߮�G�=WKm��g����y�K�&%�������#�g��F֥���7F�Nʫ]E�%Ӗ�py�MY����4@E�a��>�GV�;�f��"[N1lM��ň�;&& �� �}�Udg7%n{��D�qOI�Ꮀ�E�����˟�ɷU_d�5����]�K?>>02��V���k� ��3]3��n3�$Ԗ�� ��2�� 3�<��Ԓ�x�&ʓx-��� x$��A�b����YN#A�
�.q|�Q��n�A�7�j�8bV �}0∯&��4Ǌ��4Lŀ�Z�5�����06A.���O<�Lyv�,��T�x5���5�{��U�$��جV�c�D��W5l4A�ؠ����^��DjB�iCjM`��0"Smw�\��`���f1��}�ԫ����>��$�R@kJ�I���;���E�Ð�u٦��۪�>n�-�a����*{ӍI��7q�o$�!�q�>F��qC�7�S$��Hg��g��к��i�S�֐��.tFR��٠c&�7|_u�
��':`�ٚYU�J�xl�i��E���C���"���t"�7`��5�����j�5v �0�!�� r"�|V��O5�B�c���mf*P��S�_�7���I� ��_��=s�9�Zq���S��L���� 5Ė{3�{�nW�t��o�<Y�ĀM'4}�x@G�
�ob���K۶@�շq�W�&�z)+Q��Y���O�Vp|�m���sp1����W3=%@�"�`+�e���Aa��XlGۓ�)z��@�L����-��C��U !2����z)դ�1��������|�7�G��m��04-�����M��]wi��]S��xvW�@>�OmD�oɤX�}~)�j*�?��R��y�A��
��A�	J�	��9�S.�L�6,-+�Z�"?VY���`���l�����Q�[I4\�� �l��O$��)�=��PfR��/����J3YzIÌ���7�Yٔ�E򝒹�"����n(��H�A��/�7
bz	�����U���T�Q�)�l�C��E��J��b��ʔwf��kf�����U���T���o��y���M� �L�}��nb�é���1YD@a�U`�̷�{�ò5�Mu�[uƊ��jH~;X����[D�<LùI[T��z៻��������q,�o���K��B�m,�{��<R�g�i�S���}����5J��j5��ȿc��!Q�B�%�F-�1�UFn�2Lul�. ���Y��pW!M��Z��z�=�Rg��u2w��$�#v�EG?�n T�o�l$V�ߤ�D��d���$z�~�b����6H���o�|�g��׬}~r�$IӔ؋k�mN����F��D87����ː�_�-�����t��"a�'s~TJF�8w�U)@7ȱZ�~�$α�����]��9,[4Ha-?H?fJe��b���>��`���jE��m�cRZ�����y��s��g+jU�f~L�T�S���΅�>����j.Q8�OO�a�?/�	��� ����<[��� Z��vrAj�����ϩ�`�t�>Q@�fF>��f"� �X��N�`Iid��� ����\KĸxC�}7��a�[ʧ�W�X�񅻳'j��W�AZu�LJX%��o0G�-�� ��0���G�yo����]�vB��]RkIE�:1M�7����m�5��T6���f�D+��<�ϵ��2a�Ľ=M��ok�$(�;�B���}9\v�1˳�/8��
�Sa�P�Z�`;���-���0E�$_J���j�����R]���Kkv!���1~���@.9kO��ґ��c�#�E{l%�
��jbi>p��>�dga([����'1L	����Fa2�F�g������qSB#t�A��[�׆e:D|��f"s�%�^��<�n�y}@۪���P>��k?CSf��p<Y�����M.����Ѐ��Y�h����0f����L��@����R�X�:#m,���0M�ɫ�^Sۺ�����;� k�C���f(�$��w�-���j�j�ӝY�D�wO�en���5�:��4�߼zu��*�9���j�����a#�P�9�^5�Dq=�8|�"8F$�QP��Ҳ*�Cy��1����V"Ǜ5���;��#nO�"��.�=Q[ݕ7>�0P}^&R��|8�S��D�����]�l��C�Tru�̎^���=�f����r�,��A�)�Je4�y�Y���F��e��SF�V���"��_6EZ�t̀�?�x���Ch6���I�.�;���ďi����2��t�.Ұ{�Y�*�t��2�*�ɷ5�6��*�5�W*Ѳ:~��.97fRB��?]�,�oPyl�*������bT�^�"�E8�M����y��H�Z��њbG
՝|S�I��e�<���=h�<��!�������x��y�@��iu$�6�7
�?��5K���z�Ԉ	�}:	�\� <��|��*�z�Y�`�0���z�PE�!��7��		��s�4`��v�3bXI-�O;R��ɱ�PC��P��#����>�kJey�F�]�G�� �y�-Ą����%;oL��:�	C�Uޔ��Fg��{ۓ1֨L�~�\�5o�Ħ=�q�l��	Nts�ҷ�k�B
�F��-9��kn8)����R�͍��~�7���i^�=N{(�"�z��pi�-�,}���O��Ɖ���_�"�1�X	�q���x*=<�=4#Е#b��am�a�Y�b4@:�_B��P	�Ur��kFLN�b˟�>"ϜV0%�޾�L��YJ�=��Q$�F����*����4md8N�q-�/�}�>^ի���[ ����@j���D����_*�
b���J@�׌��u�\e�<�e8mg�h-�K��:7R�g5&��d��������Lˌ*�;��F����Y���3���^��M��7�:Ž�&�]��B$�	�	�d��Aɹ^���Vyt1{<��y�-�	�)�� ˑ�#�?����@J����!�4k_���n�%�^\e���4���e�:p�L\����X�sܼ�2K6�?M(#*���g�Fϼ���%Jpt+Y��Ӕ����\�[	�bg+����\yӫH}�	n�R{__N��X&hB֋��g�"�@�����2y"�v'���It���/}8��"�C���@�>X ����&O����\6���Q/��7c��]'�[�/0��,R����ٕ9�o��x^��U�M��ו�I�g3���wߟy긋�i�i4D���%W�m/g��/dy�/�V0�8*<�-匉��~�
Қ�X������\�#�����8{`�U86V�{$������*�ީ��E!�b�!�D��7${���s����h	���O%}'�?�� �z{U_pk�S�-���ܱ�+�~��2ff���D�6p�CR-�բ�G�
\|Gȣ"�T�x����1Z���u����Y':]؅��9��K�p\���B�ja���?R= ��t��ڟ�ެ�2�� ��>xN��T�5I�b�p�iM���H�F�D��?:����
���_Ǥ�@C4y����]���@��;�U�RS1G�uT�Lq�H���rT�V�D��ڨ�坵�'�J�%T��M[p�D��^J�{b'c�jB��:���P��MB�E����Tr����`*�Q+znڼ���R��1�F=rDGYk��6����a�!u���D�|I���"�Ɓ䡔�ι۱���� ��<�� �i���r�ƞ��N
_d�����1X�Դġ��F��l��m�V
��s=7����T�.itۂg���)/�䪠;��(̗H�Y7ݖ��a���y�n/�x� ���z���n�ڤq�O�9��!%Go��L�
'�,��	�<�4��v}��i����A�ޏ+r�Ŵ�m�՞�;q�K�m[���Z���B	q��[�C�m��A�뜅����Â:�洑�fr
�/څMA����m�QdE�_9�:�jM�ns���nb+T���z�A�G��A{�I�YkR���л�d�����Ϯ��?��d���5,Ӊ�ȡ����C߯�K�6���9h뤵'��UR�C,�5e�eǜ`x4Q��^M�b�tjW���Y��{��o�^��3>$�%/ӄ���Y��ɽ�-í�I��C{����oW��:��)�D3R���$8��s�:���}~�v�G1.�:����s�V�&
�g9v/\�S¸�.W���\U�ޮ:I�(��ez/��.�	���x=L�>��,�,�����Qoi(]ڿ����|ec�>�N� � �BO܆_�yAT� xtC��c2W���떧O���i�}��� `CUQ���4\>Vh��1�T���R�kjцs]J���N�@���is�\j��Eb!�?F�<�f�c�P��-x����8܈��8 bA���-e����A\P�����h���g��5rO���T�`iEL$�S��ه���uJdײa�|����X�1,a/Yd�L�4qx{�N#}e;X�5�15�g���Ku���0It5�2�R�{-�v-}�����_�y9i���@�3BNZ���9K���8��pYe��RHi��r3<�������\��e�6�F�k�x��$����Sv��D��[������}QΤm.��c:�Qp0�~<�L�I	��bQ䈽R����#ap�{T��lt�c#���ƾ�y����#��W@�F/�^��`�X	6��cT�=%So���J~�uI&����+mc���;��]5���ו��.K[��)n
%�c�#i#�Ivx"{���%�[��#�9���/p ��q'�a��D]�/�9\f�u�!1U�@\��Wu�2è��!�c�<��������)[$�g�|{#6�m���l�`���(��� �̧0'Q]�!��aU��m�9~ĮLzՆ��h���N�`��+��t������ǁ4�?e�6��(#��\2:L)Id���?qe��R�D8c�J6�{�g�~$�Nq��S��l��T��ޔ�{����ȁo�}�A[�`6ZF�Q�h`�M�2�2*�F
���c$\	K|�%h�-DI0��R����D�`k�_��=c�
D�L��5A? �,9�
D��M}R�dsWF��ᖀuAw���r�
�RŐ��k�����b2\��������i�]�I���JQ�ۘ�hn�u6_�h@��ę@C���"(�5�|H?�<h���5��ou�'����m�%��t��V ?c�P�Ά��va�ʃf�x�0`�Ȓd�S�p�a���/X���!�n�:F6$�|_�QB�1i�@��(��}��h1薿�$�d���sk�\r�ӌ�r�"M8IT>�?&f�A/C!o���ŉ�L�&�v=�`!T�"^n<�����/���Qi�~\04q�j�'�Q:����6�ծ���l��<������N�K�Ԛ�pȸ��ǽ��=��_������d�d��踜 ?���+x����LBE
	,�(�Q���TZ�q�Qq��2]\�K�Ep�� �Oi
���0�ԯl�w-КF$ok~�� �j]ȹE�Zƍ�Ē\2�<x(mZ��Q�]?���ϯn���^2�૫��)��?z0z)R#~�����&��1��)
���B��+�Zl� �P��5���z�;��͚vPQ��#e�=����zV�!yff3Ezǭ�ܥ�ؑRt��$,��ô��l�=(�n\{��e��K��+v#��-Ps�)e�t �uGw=�8v�h�و���)��[+�G��.Y?U��%��8;-��3O��XR��
�s�0LSW�lǏ���"�E*s�a	�[�&�Q�88��d�]Qm�j"�j^%�� ��g�Á&�vF��]X�6F��^�֞�օ$�O��j�EM���60�=�K*#̞o;�~�46{<ƭ[R]�'�Ԅ0��/?r�G�t����q+�2���~�M^Z�=q.��'w����)O\��I{@<[g��
o��R���"���7ϲeߨ�j��0�qJ�
�G�'+��t׸��v�q*�~�Y�C����(͔��&���S�cu���e-49�{�܋T��Z� J���jj��u��>A3�n9��]�8]�7�7���X%!4q�5ԅ���\��ⷘș{��t�� ׈t</�ȈБQJ^p��� s��%�	��qeiZ?Ժ��q�O%�%<>�"o�þ�֣A�:�{]+"( ��������Ꮠ�)��/�{�qS�A쿊St���{�
&lma�������	/�E�ʖ{F�$������4����6,��b�-C��q�J�o��N~�Lëk��S�N�QI�`��������w ��(��u�Ȃ��_��$c2E��Jz�p��~������N5�]!�{���z���m�T g�(�����=����и�Fd]^gֺ�s�i��'�<-�nu#���j�B0n�j}f!a)��/��u�_�':�$na!�!O�N?���9���3ڶO'�(�A�F�?A5�=��'���TÇL����u���V:1\)��K\��خ~+X:W��6�h�`��c�7��P��3^�\|�xF��3�o��!��/^6\�����_�Q%��R�	?��҉ջz�IP��V3����o��wgcڕ\;���V�/ݚO��B]�ŉ<BsgI��3r�m@���]i x��WL���L�1�p3��Un͵���R<ki����,��IB�� �G��������ap��2w��;�j�+[��
Ѓ	���yM�T�
�u5�i��*��TO(��	������7b�j�9\��CSϕt�8F�߸e�(Uӛ�3����q��Z�Sߟs*
��Y�Hbx����(ӎ��'�6^�rʼ��Z��o.��lj%,T�G����e����t%vV-�-��IqmK����*�9���C��p�`�S.�4��$W`L�x�;�2�%*H�K��R�"CEac��)T��s]� >?ل�_���������֝%+����$<D.��K?3j�P����m���e��55��,A){|h1Az�F�]�m }�W��l���W��"(�3����SȺI��	y_���g��|�0"7N���^R|���^�Y;��'���X7�bX�)�9��K�{� SbH�=����U
EJ��%L|c��Hth�f�A��E�1;EQ������e����2�?�)�����	���W�'T�LB�Ax]�	�`��5@��kC:U�z(<�	�x�5�O���ط9-tVX�hD��W�ЮZj��\q����
ҍ�A(#�'�!Á�ç~�6�,�I� �ywf t{5[&���+��r�޹F���u��]������r��Q쩧�XFό�����giJ]x\����I����7w���%����ZЅ���Z!O�g��ą�z�PG��Yk�!�=dzrº��C��~L)��d)M�<�����<"o�]~��:��z��
N�IE+�c�r�,����o줱���6v�D�W��{!�R��X6�N�B(-��m������(�y&�3\�T��0|7��^�d*ԩ�!\|G��5Y�E2���f�b�h�j�f�n��y2�>�O���.\� 	��L��{sL�w���#�M+ljJx�jt��yq�Ľ�LjP����`�����G3�_�T�a�.�~y"�>^Q
�ïߞ�M�4M�ax<�f��@2oC��CQu�G(����MF�a��d|EH����0����`و{��*���|���{�C�}AR٬�i���̰GnLg5�5�
�d��dVց֟�lr
:��AkV�&̯��yRuBձ�mW8SВ�Q�݂���P�2�`)��4n���������b={Q�6��r������48�G_~������b^�KzZ5	���O�*�v=F�7ۢ�w烈
ȁ�g/��d��+.�f
���ڕ.�3#Q�0/
��MO����+Jn c˜��-�<��E�c��&�`@��k��������8vi�e�v�+�����G���PP~�۪�������UBf[�C{#�.���al@�;	I�?�BR-/3�`d���E��^9��Nc�ap[u��U�S����Dx��=Y��Q�ۓ����  ��CQ���T��:���{?�(x��ԏH��Ϡ�d�<��:0�/���飫�G�Cp�6��jW�!kw�0p��;j�]�2�`��]ב�1��k����C\=���m��h�r�8˲�󝿍�~&���*D7����ҩ
���ZwT���@�Wc�R�X4䳼�ͺ�=�A�eJ-�\�P**T���H�W��Xu|qi��y����f���q���390�%����.����3{HtoLl������j��r�e:�1�^�8M\)��:���T���W⨔+�e�eew��X�ˑ��l�<k�T,�"��uw��RV9��h.:x�\�|���Ӎ���@X�-�=���t��G�H���A!hD�������;���bY"lm�;�iW5�yN6�U�`d���?B)oE���&!��
1��U���Z�m�5ot��A7�k6<�3�8�v�E���o��j�׏2���kO~�>4��K9S���Z���=� ����	@�$r͐���ו���~�8���n6�K�_8/�Ie2��qZ��߹ny��X@б���(�3tM� �n'LpJJ,27���T�Q~���'X���HD�Ψ���a���m-�%�&DA �����'��r�����[��W幡���6v~�0|ҡ��"�'+����c+Y?έU|p�x=/s������2 ��Gv(�ǘ�b��3��ށ�n��.1�PȥX�ї����v/�����Ʀ�Ex[D�o��>tf�Zf.T�yL+��v�V����[���Q<�0�$�1�뜺ڕ�n��򹙝TX.G��
���^��j�4kq́b?š��X\`�u33:��Q��ڦ�S/l�Ɛ��ӘDf[�������v��Hj!ݢf���.)yX��_��\Mq��H�~>j�Et�́\���I�.����ٛ]E�2._�x��Y��{�R �W�i�&��x���&G�o+;8��!/N�Y	��ks�-����{�rx'�N��y�S�mv,�t����]�;��)�k]3]�F}�n�e�	`�޶
q*��)��u�&�y=Px��-�O�;#�q���)�MB4�(1�)�.���vZ댫I+�o���� x�wzFbcE4r��xֆ���I��[�`7��X��5cd�(8�3�"[:��:̏@^�el6� 9�#�/<�U�nc��VXZ@�kң�����M{����FsOx�GbU~�sGJl������֓#��Yy"���@��!�><9}���@�a��ܺ��c/V����$�lt ����,��,afu,���Fm��)�W���w�x��<;If����o	��G�΃9So�힩w�5$0�m�J&�J���<��^��������n�kG���~����-�
�w%n.
��
�$��G 5i�KI��j%��3\p�7d�J��e
��j����wH먯��Y���(�yQ�:h�ۖ�3��Ť������,��{L�NJq>�C�m�t�iSi�����;���pQv�i$��r;�E+�j>��7���L�}qQ�O����f�Tc&���1ɚu��X9��!n�?,x�����"CB�������Qh�f�{!���|���o���Ն?[)�jEWd��Rʖ�)�.9%�k�?�=}�����qX���:����%�[�����f3d�;l��컬d'%�סBR�T�F��ł=��d����-��*������졄^N;d޵�JL%�B҆�n��9������U[Pa�OiuX���-�Fai,�*b�YI!p�p�1R,�e9V.x�+�.G�65
�����!˿�Y=L�F�Š.�+���U3���7�9�k֎��Z�L{�d����S��q�l�@#bvv�M�s`��g����`��D���Z^����0��������Tw̘'���CnzY���@�H2ogܻ�X�1!=��/�\�+/5��sEwq&�-����r�t�w��� +4�� [���ޮ�����@7 �{^Z�t���F@#n�;9�=,N!���*Y2��ݛ$5r��X�T�l��d*KL��I�M�zU��:�Pt�2�e�]&t�O��ja��b����"� ��|��NP;�Wp�Jچ���1A�.�R���T�,?v&���޿�/؍�SA�*`s�Pz��� ���Xm�˫�:������+K�����a@�*���n�BA�m,00*��8�9���ny:s�:��c���] I�Lѭ�.j�-�%���3R�õ�����߭���ĭər
:��<�0�B�O������%�S���rR��*�u�S��4����K��'�{I�#$�{ns�n ��3 �ۂLRX9�P@�ҁ��h�~0�/m�m�}���N?��G�����<Lב��ؐOR��o�R�<JBZ�frXee�vʹ�l��%�Ԭ�*u^�k6Z+;�\$N\��a�)�&V��7de���S$�9 dEu:�ȁQ|������HI������h�WgS�<�CT�l7�c�����OT�T�:�f:�ggI[BZj�=��l�2}�#buq��۸��?��G�������`j��?A��3��_O�Х��-4���Q�y]?����@m��3�j��f=��ج"s�'C�^�V��怩��Ǹ
��Ř7	���AV�J2��4�X5=��[�n=AS��יo��~U�&� a�9��1���i[�b�{h?�Xta�����b�RN7��e��\:�X��-��+�Ԇ2�G{�^s[���k���E)H�N	}��sEG��J�U�ճ\������/�i���lc]C�`\��?`��Ļ��Q����\5(���Z棺�ڻP1�Ν��Iv�۝��C�qt�������0�_MBw���R���-R۩�eQv��lH���(9��p�L�	!ֶD׶b��)��*i����˪j͟Ya;9����"�����v�e���a�����~��\�_���TF����N�L c��o��-�3���V���.Q�Bq�Pi=&��H�'���{��J�Yc֑޴�i6��ܾ�ib��0�l�����i!�"����SZ�%C��$r�@[R'�6B�lb����}K`�q�i�-�� -���k)*G&�}��<�GSKYLh��t��	�y�˜�F�v�kz�q
+v8j7���c�ٙ-fCP�w����#����F	�!����v��5����	H��� !,���yL��.�@;�+�/aG�jy_E��%+V8~���0��F���
��.�����A([���'�#ƕ��x�O|�^��X�j�V���ZW"J��V�$�BW.���g1�G.�����7VfKd���K����"׉oN�%������s�6	�f��5��{�<�
�����١k��l�� ��������l�:��eL ԺA+��#ȓ�U���X�Hc����ˉW8�rcņcAn5Kb�w".�:U$�Y�}uO�l��M*�/�{�.�����K��
��j�"����ڊ#�sQ����ȸ|:v��N]4M���[Ӑ��8��(��T�kґ��[/�z%jCd�z�	��u�g�����������[J����#�R�Y�?�1�Ѥ	Q�j�4����~R�*4�,��������8DE:ı�ī�b}��.����Ĳ(�����1E�qlU�6	Z3���W�h�@NiƢ��S�@�mʫ��G��/@�)���E=��8�K������O��J�u,U�ʹz���b~����Ī�k�T=`#���U���������f�3�4�پvqT�6B���R�c�:��+\� -���	��b��'XM��P���1.Ӏ��X�����$u�j�G�d���y�������X�J�h�t��5�1�0�����X�o�88+�{��/�xv���x_N�����m�L2��%�h/�1�%s��|�=
 �1�͔�o"�tvš���º����@�e�B(���PE�/U0$��B��b�'I3�
���)���i� ���.�~��L\Gk�$ �b]d0U)�3V/�p��$�l�c|�i��Ҷ-QY����'�L���ð�U�����JR�F^��?ꁁ�d�R�Y�G��u�%���|ȢKHop�U
5����~�z����3U_Ȅ�Z����5��g�0��ª�����V׋��y�:�Ɣ�����?���~�bP:�x���(���aQ˚��o�㣕� ��%_�*_\z�����j��3�����$�R��z8��0��'��-q�=#�7k2)�s�1>(_�vAm�Sob6�݂1.;��U4���ÉDe^�8���y���6�y���Vzs���)����v����$�`q.�WbT~�4�H
@3Ś�G��ǻ�<�PWc8��>�j����yQɝP�!���Պ1;Q?q�P���k���+D�4�\y� b	I� �1>�+ɧ�*�Y�E� �.#��gU��j돇� e  Ϟq�ܺ�(�0\�W=�y29Gu8VΞ�4�rS����[T�Oo}����H��g�];����%�h��6_Y����4�#�E����ɮ�y�� c;���W~ZP��岽����LN�1�M=�{���
�۝���c_3���#v�p{��t@�R��V&7�*8m9^�O�oói�k��T�?�6�#��_��s�gP!^-g+�o�ޮ�[�j1!>��칖j�A>�~pE�+�����8��=��^�cxp�Ʃ*k_�0wj3x�_)m��<`TU�L`��QJ�����?�)�9�W�n��	��ί%�%���!L�Ͽ���<E��6yp|��&XI���U��ܴ�t����I"?W�L�w�����ӗ"�������ɿ����Hd�|$�k_�6�0		r�0��3�I���ǎ��9�<D2�|��6k��H����'U�9 �(1] t>������y'c��V,#��J`����܉P� ���hb��ҡx]�1X~�M�h�K�p���D��9nt�>�禚aܾ�f�ݶ�_H%�[drL�V8��@�A��~�� ԃ�:�H��ݵ^��}5���a#��B_��H�tP��ۗ�t��wA1x��l�k�������u�U����(1|�q���]B'P *����kt�j�ǋZ--�8��m�$�N ^�ۡ�<IS��v��>d��@�w�t�f���u�d��gm{	̍��B�M�["C��΋�_�\����`������������:��j3M�﫠���M0F(����w�S+��4��<�qGul3�Z�_��@	~�1Owc$^��2=�jl�w�{%?5\������@����)Ώq^��L�����5��*@�m�I��g�
#��
�>�a�2�r�t3�<x�ULn�g�8t2�k���5����W�a�G9H�p~�I�fї7�q�\>v*��=*��
�>_���F�V�分1Gl'" �7�����ld�'�P�-��Tb�\W�sZ���wr��,o���'���y^�u��>vԀo�I��S��h����u���O	e^���Y�Z�Q�(�	p��,-�D�l;��I�\��"'f��&����Z��9��@��hr��F�iA��)o�O	�ە�l҈c����w�}�"�O�\�8C��ˈ��q(�Eh�P��ک]�W�
�@���)+`3b��_�wiXI�)�{�ڶ��Yr3�gV����,���%d6	�.�,��U+�����6N��C��<BjD|f�0��i֗�{��1�v���6����<�Nj�%̧:�ζ��k��d���&���3�Ä�f����H(����>�al,^
�\}�ڿ5���l���y�[#DX
ޱ�H@qaY�E�n�2xh&�p�/���pZ�����]7Q?_X
)"yY��˿88�^h�8�=G]���+vw�~��0Uq����(2�ӡ%̂FHM`5�O�f�4���@��Q٨H�;ǑT��=��<�o��v I\�C���>=�o`}�f�/'�&"M_�3ci�ז��Y�5�/�ΕKXs=d�k�3���?`h<R���ŎZ��S{8����Ÿ�|� o�CD�m�Q�A� ��VȭR8λ΋������ ��Dde}XP�c�~�����ePH%1s�Y����%��F"�;��/-7�3��Bз���@�~Q��HL�?L��v]��>�l��?
+���bz6�u�{7�+ǝ�]G\��#�6���b1ߙc���4��	J��N�No��}��@�:�Ų��	[���[�%|;�le�9��p`+��_��$�������-�����n�k�\��c�9l�����j��?:/��WN.j�N��í��s����u��z�����Q��'D�&w�`�$:��u�t�@�^bu��`E�+��A�A�N��0�:C� �/.�q�_��_X�f����R��,7^૷lV���X�1_�#�z~��Eq%������K�$co�c���E�
�C��u���ۤL�s���TN~FwT!�,5��1%��8�M����[��D/��܀��C-J�J��-���Ab��������5�E�MC��Td0/1P�� ׽�T�ݢ
���/"����Tnµ�`s�l}b�"dvB5S���[�Z*Hv�����1����~�ٞ����%�+|*���q���m�7d�ă�a�4Ly&�pVp�s奏qC�؞֬�14C�ؖۚ�FTi�ib���Iy9~��n sB G6i������'K�V],n�J�^a����4-�H��zB���}�`xV��z��ሀ�׏���W���3`qr�)��"ؒ�o)��U/�k�9���e�<K�D"E�'��jU���8��!�
�
��� $�z�4[پ�?Qlc�]@����?������`�|�����8`Y~UMJNOH,*��C�rU*b֊�#B6�ͤ��� ږ���e�;DSX�x��>{��i��b#�=�K�Y�g�߰�����j��۪Z����*�Kɋ���E�cgG�����ʉ{�?� X1Ǌ���]E��KOoг�o����� י�~z�´���$�#J	s�E�]/~�Y{�k�>gB���$�fq�Y�=��i��6ǰ�N��D�"�s�/��1�+x5�=O�� 9	>:���������b8�P״�pR���C�ˬ�6�`3M���Е�Fv���Tլ間���&\�����Q1��{\��֗n:�>�_Z�WW,��$l��GD����l���ɳ3��y_]�����k-��Ѝ^���Spk�8�9h�X�4K����U>�a�QT�W���U�?�%����r�V��j��1o�& �T}�}ou?���R���
��Un���mu�=|z���Q�{;���;��Wea ��4VB��_SIL�Su�zH�(�Ll�g���grOV��ʝ��ѫeK9d�ګ����u���"*�Gm�K���|���;DNL��M�8��5~�F�GA��_��)�����حK�A'Ԕ[�vݔm�H]��7N-,�,P�=���J/z�a���>2�����Ʈ�_�'n�n1���I Pc�Wz11��W(�*b3��2F��n9O�H��F/����rH�Ei&�.�@V�J��s�'�J��&
%���T���q�&�]JA���O��p)g)���+�#>��N�~?�gT��]D�1��[	��Y��Bg�u�5��:0j�5җ�u�m��y��l���d1Ovvh��'��:�!GQ=2.
1��%�@ݭ\�3���eB�X���f���]���W6�a3*�aerBP^����z��ƃ'E*)=ηH���-�p���n;��b�;:����6

y>+%�����o>���c�z??��N ��<��nVPhK�qƚZ�К�ZeTI��4�W�\�A�-�=E��R��}���(,r�u�(^H�$\�q������ш�`2��ȥ�w�
x�,�Vwۡ��JP���2��2d�R�J6õV�Y5
����2�n�626	��;Ng����UX����\ۍpF;�Mh��z���~۝��F�Y�Rg/�RX��V",��N+?��w��k��1+X�M�	�j�G;�s�)h{���͎�o@��v��Uyј=��@��;��T����c�*�i ���h~t����Y�;p�*Lw�y	��k���TYc���u96���	m��A�<����cx�_m̤F����C��*�QM���6��`��ŋ/$�k�-�_��7!��&���}��f:����˿���"�a��E�q����i���^��X9����0��Z78��Hf�,�wq+���}_�~�;�����>|�>Յ���Yḽ�;m�?�$����������xr��lאGU��bo?4\�Մ�6W{j�'���QR���ǐ3�"��]%R_+�J�g@yQ�� i�
��^ɑ��	V�<��8��M
����&/��H(��!'�\c������>��KD裝�������	tf�Ͳ�E���?`��O2���R"ٳ���G5F������?T�Q�� �J���f��Ll�Z��׺:l���IA�K&-M��M�,���+��i��5�Pݓ�*�^������L��Xt��%���DDV�s��
4@!�p��^�U�q*%�{��s���.���ަXI��'�N�y��=�2Ò4h�n��	��r&���zs�^؟D}���t�R��`ŉ�O ����s����PU��y��"K �:�'��nU� ��B���.3Gc����_��)~YM�e���\%����3����v$�$�%�7�5�fI�\5%uS���:"����]�L�9��ٵ"�2�-��d�
����RP��(�~OW1�;9�1�׻W�����th�\4?�tP�y̌r�N0�%��`��4����V9I�  �/K��:+���?A�2�OH���;�y��+3��[G!�^�E�
�_)n�'�j�LtY�6�YY����s%���ھ{�H5�w˰�Ü~ߩ�G��|���I�{3{�cIyA�S��l9�4zJ�~q���<�9\k0�
=�������=��iV��< �)k2z��������A� �lE�r�����19N��©Y����?�0���ķ�f�,�,{v0D�,��C�̧-��Z:]�^A�e�=���q����,��������!o����=��~�l��g'V����)�'FQ) �v�Ƒ@��C~w����w�k(�Ha}���]��ʆAޱ�S��4�vi�9����;Ҋ��)7�e��� 	�
.R���qr�^��6�ϡy��u;\.�l����^#@�n�Xn���|뙤�R3g�<������8��`o��v��n�H3���Ov�;�������y�φD��X�heb�^സP)�sL*��Ji�<&��H;���meml���	��OQ�|d��]�/�W}�zDr_`����\�*K'�j%�t�����}��+(��v~d��@��G�p6ݖB��뫁c��l���G"���]�����GJ��Ĳ�7�G,J�4ӓ-��U��$�_�.ܳfb2�B���(��;>�R}`
�I�jY���4�:k ҚTI2��)X��K4L��p垤��Y��T�����L�*��N�J2�K�M��;h��l�O����i	2 4s�^m���Lc�L4R�B�	@]J���{�Jʹ��Ed�-~�چJ�@߶��൨���L*0׋��a�>O��rj�H3�PJ:�1i� ө���db�������A���\�,ܾ�"W�!g~߸~�b��҄ǁ��Y��Ǽ���+�6���r�E	�I~��kL��u��q�t��s��>��_��-��!Բ��@�K�l��w��%捘��,׺�?�ؕR�Ee�u���R� Cdjf��9�`H�!aЎhH��RYT��*�W��nsW\���qna-��O��}u���Jo"�f�d����Id��E+��\I�Mu�wl�c~��=�ɦS(74>�ߵߩ� �+Iϱ<Ě���
���cz8�0*�� �$�R/e�/Vnd���.���r��dwP�L��(o�늼�[v��=���eO[��k��<9g�/�Ŗ�3 �ֵ����U���~�ж0�7��)���ߝ��:;��Q}�DI����1�����n��hY���2�-����\\�����hx��e^�-C�*�f���o���zT+q�/y�����Zv�a�����3R2-v�����;)Y���z�v��)cs�T�H���e�K��[��9�1و�E\`��	�u5b�{����)�\��v���E6�F}�ذ�W�*m��ʒM�	�e��N�T�e�hjc1�����P�6�0���B ��)�������|�f�q,��J&=���i<2��<qE=PsV!D���f�Ա��0��anQ���-�K�2��R~t��F�Lz^�
�PxV�u�7���9�g{��'/c�$�;$�:ޅ�����-zQ�����E� 
�a���bHyEa9<�Eh����;��|�l�60�fV��t�?s��b2=�:O���x,pZE��甪)�	Ae|�T��W3<U�C::$��[o���@x�\�z84�I^TY'$�5�B>�x|;��iE����fG,
h�˵Ӗ�_E���Xܿ�v|q�3
���䲵5~�Q�`�����|��5c;:����8H�YIh�v�o����6*�	ҵz��U)kk<wU!`o���s���wě�7���v�i��0ŵ�����[��XJ�;Մ:�.�%��kƓ�	���&ja_:�1�q�J3����@�޽4�Ԝ����0!��4�ᦋ��Q����YՃ�B�����j���/E�V>w�����.�GY��j�+�!q^�`��<9���H&ǓR��Ǚ8~�U��dΘ(��u�	^���	K� /�pb���0���%��>&�_�˱ !��]��������,�}Fh��.g�
}c�!5���_�ʈf+�J��:�1���u��G��-5�D���)�JF��ˡ��5Bb���
c��gQ�Up�yGy[��E��������m��74�G��R�)�`;��<z-����2�%ȸ�@�.X���4���S��ģ, PF�~�j��Q�[Z�:y�ibfN��+��F�-X��h�;>лT�q��m��,X$�l���N\1�)Q]s���F��z��
h��p���ɂ�ց�3����B){��K9	�hj+͛��]8��d��!f��ϱ�s�ʦk�ƥr���	�z #�4�ڼc���ĺ�L)����Q��@�*Q�O.�g���������V�@J�T�ưX�S�d	�[��\�U~X��l.�id��� �92b���T�[���7�7�}���յ�w��v�ei���X��%�^*��"��������b�/O�'Tp+W��2�	�A��M���)��n�Ю9(�<5U,�x��GcP���Iӊ�&IK�\�.,������*m�~&ep�c�M�o^?���#B�U��B�Q#X���RLsq�N,UYJG�$Y�!.ޭ-�
�̟�B6.g���`�`�V�*��4�<�����0���~4�oY�!��ml���/�'qVLF���|j�V����� 9�r���5%��W�'�1-�9�<r�n��O Y��4��~���>usSpR�%���ՠ�f�XG18��O�-����#?���>��k��/���.�6�+n�@��VEV?4ݏ��K����O�]n�1�i�����£sE�Y�c��1��B�� ����C#'���pV6�,/~��A���@>s���`�rs���$��ҳ�$�H+����at�,�Ӧ9�A�j�)�r�`oKr$j�9�07� �R�.AI
��T�/�3-�	��+~ع�$�64#h�y��u��^^1`�S���O�E��
���-�r�ǛhT���B��Vo�
1�a���X)�EG3��|����/��zUO���S��5q�*�ٴ�\$u�HL܏QcE�Q�cn����<�w#���R��b��/�a�h���'�/9�^��p���lˈR�,~ۻ��O����]�S����}�-��t���Н�'M�MPv`���B��{(@�X0�UK�����.���w\���X�X�C�=��� �E��k��(D�$59)5�7�~�hИ�4�>{t������$�ߪ\�q��bz�`�3��8�w�ޝ�Y)O�m|��&c���?N8� �	�v���z�s>z�.Q�[n��
���f��u�����}����tk���d����js�#�u6�/ۊ�~0&yL�6`?�Y/U5����s�kQ� K��ԥ�t8�aQQ:/��P���t��.�l�o<�K<(�#8�^�V��t�I������ �}���oc90��=�Grt�L�ER}��|/������2��L��]Ѩo��^+�?��)u�Y�J�|�t�y��`���2~�K��~� #m\��ev�}���΄��O@fY] m&J�!tޱ"�X�ޕΈ3Xr��˛����e<d��1�r��4�$�͢Z�"0�~�q���H�R�D<�u>�P7HS�)��)�䠼�W�S �I������M�B!�(�.�6��:H�L�C�[JXy���)ӻ%�+�_�Ur܀UGrE�y�}-QL�Z�C?���{��h�����_���)I��3�}��j!r��N]����Ic�
�jJ!v伾��1�����Bs{E�����z�t��?R�����nTls�Ṇ���Wz�V>�P��mW>��+�:�<���/=k^����C3�,��
m����<}Ѝ��nTxy�� �
�9���'c���nG��A
���[5�4C������R���_
7�$Ra?���z��( n;�XچRӆ�����8������:��&Hk�L���`��G_ѯ˺R�!T>-�����8��sڏ#�b׿`P�@)./�1i����,��������;�)��@��M�]3��	e\��l5��ql��qtu&��5��+�^^W�}m�z{��Z!�m�H.F�*&U��bpQu�4x��_�ɐ��m��ȹ��XrH0��v�E�=�E�b*��*�a�iD����Q�����f,ٌx��*��r���d|�r��b4�w g��gG�8��1X��%�6�'�J�����|e�o���<}4��R�<r I��`��V}W�H]�=�M��*��u|�� AT���ܖAͥ��R�UEH�2:�B��ɔa�<��!�ػ�t,�iOve�k�=����QY��6-r�J�����TM۬5nԀK;F@=�]r��nR�/�#�B�T&:̂�e��ܗ�ׁ��Q&�1B�XR.a|%>�;�T�9Z�_DӘ�sk�����GU�����K :��:�?d˅���(��,����	.�(�\��(�X��?�Ə�Y�)�/Ԧe��_�&H�7x�A�s�he	�0�'q�Gx��[=�2r�|�t�1����DU��,嫶S�/���/*�23a�]7�Ԯj��em�xٵ�H�ќ�V��:�ȆT�N�`����+��{M3�_�w� Д4��C
'^T&�c�PX�|4�f�^����/�ey���_>&�[ʱ!��M�;��0��L�{��{&� ��؟�u��d�4c��0#�FX�K�Ki�KY�b�6�Q2qv<���������)�md�-Hz��:�$�j�lbit�!��u����e��[�Q53�l��©fB��8���ю,f���Y�X7V�轴Zn۞ޅ��?����V��M��.�7��&�aɞ� m1�W�ޟ� �B��a[�х[����f�����^�h��G��wn^���F��6k�B#��u�G���ᕃ*�-(P,CR�-����xꏰ�Y�+U܄=�*]��f�E6�l���]r\ɅO�N)X��1��Q�
�7+L�MH��&Q�n�}���gj�Ya�^ا1�z�������yqd�_3eY;�y�1DH���~|	�!�\�Ѓ����)4&��.g����ʂ�)������5�ϑC�>�W	"��g��Ae�r؛!��ؿ����������{N{/n�82�xG��)8�ĩMMI��4���*Ֆ���`��Kx�s�d�;�*i����pJ��|����\>ũ��Xmп��.���1��[V�_:ѽ3'���Y�5Wk ��y4�YA��\�x�.���ex�����<�}d��f2�f$�Y��7P >i�bu�Ia���Q��p�/"D��p,��o@Clw�:��X�%���4Ə\��	`��� =���{j`b�^��F�V����6����]V�L	���4"@T�oaF�s�f[e�|P~��h�؄*�+!(������ba��j��2
����3%���V:L� ��	w�`ZѸUA�ޱ��Ɛ����狸
���ZC�����>Ҝ�!~98��u��/$�#�v	ε��0�}��B:x�cD��\3���I�u�
�sN~�N����,�D�e��	����ǜ(Ό�C6�I�{%�]��$�ǔ��	W�K��M�\##|�����H�Iq6��mY����w�o�r��Kc����r#�tɼT�I5rk,��c\�2��z�w�s�Z���p�i�s�6h����~�à��o�Z'LY��Ԯ��#��覱������&�+T�$`D��N����"z�1�1:?��.�pV��~{:����jt��Q�B�����C��vWK˭]�a$�v��e��j�|������*�oC�Q��}^��}�B�)'��Ojx\����
���Yv:-��
�(��{���2����hw�s[pu��8.�O3��K�f��3��Q��*gM]���!�n�ɝ����1U���f.Eر��Q�0t�v��8�z �b���N!脽���� /���Q���Yh�Y�:�vn�
9eD�Dfs���*����͑�|	���A F�������H�C��8��(%-�$V�Q^-���D;1��n��0�)�I��9�2�<���}*h�����:���<�P��L�!�ȣ���*���c�����8NU:���.B{�g�O`��?�@[�=⌯�.�o�M%�y��� i�����V�w0��U�-��;|�E��{+����4E٘���ԏ�)k:^�놣��`j��I�`�f�\=��9�3!/�	#��-��_�G�1�Q��e��c�%�~�1j�mFpA��਒��r���"���Vʥ���k�Ʈ׊f��Y漑���[�u�S�Z�|�}�K�	��&�PG�s�9�ql�u�;rZ���$xK��z������a�����X�瞁#jy��Hb�� 7��p|�ȿ��X7[ں��豏��S�BC"����?x̬~9��5��M>ݼ.<R��GRcɼ���}���G��7&�nU�rh�6C2ӛ�ą&J��3-��^HiI^�_��zt��IA=4%��s���s���"���C�~��"Թ��	�S��\>L 8JSE��:���l���{������>3Q�x�����mAp]v�1������ S�F�'�;e���My�W�BX'8M�}��ܐ�������i!��Q޶H�5/t�� �\5�a�����Q���M���ò���~��a�C�U���Y6b���Z5�K0���= �F�H��:"�FLG8�+S}"H��Bk�Uf3�Z��YD��脘���H(������#Ի��d�P��z�_sKq�B�v�0�[h��'Y�`s:�=���h�:�ہ���e'Hԝ�o)'��C���=�^�q�\��e�]Ͼ$�Li��?�:�T� �!QP4��[���G3[���S��9���yŰ*A���x]�g@�����m�R�#��[���<�d�)y�	cL`���7�� ϲl[l�^�v"$ۛ�������ة��yV�N�k��ܻ�B4.�����&����
���W��m�첶+'r�8�&C����il�*�_��X���(�3Yk��*%�Gؙ�򇋨$Ӥ��:��/���+iY�'�Ň0���Ʉ|����}�N�WM� ���^�����
0��c������"Jh�wV�b<��t���![Eٟ^q���H�Y躧U`	��-;J��/1��[ٜ.��+�8��;��9����
E����:�bzZU�ns\��|6��5X�Ba��C��8ƈ~���T�V^�b��s��j�2�0u__���/5��/J�	�8�@g��6�vKĸ��,��P���ƚF�Z	�����``�.~t�����ª
;��(Xb�/�I�ĒS�fZm�����d���04J7a)S�T�����:p�㉫s.n5���4ɔ�S��z\x��=Tg����U���ä���I�MG�#��L|.@g���z?�O���g�OY�l�[��rp�qR�h\�̩,m�Ğ�x+]�7�m�U|�9��n�x1�%8
�<�vsg4Qe�D���x�~�9l1[C�N�*Q�4����t4�� i嗣̩ �+%p��u�VZ�s(9�C����Nvg���z�T���B���xA�L;��0�!0l���n��PQ�o��B�����uv>Ω�&�̫fw��<`^�~{݅��i����`��=:�R�jY�~|A�φ�w��BY�c���j����s��=�`j�=r\q��-=��U�Kk]�c�*�6b}� ��d[���G�&L��P��b�uO�g#M�,.9���I�!�����Oa�Bvj#(��t�˺�I�$ \��U�iu��t6��0mŹ]��6�5�q�`$q���M+0��A���C#f�18s�o��_]��g63b�6��6�0�S�`��mV	�,�k�~��F��^W�"e�5:\�W���\ڦZ�^J�i�8��q�� n�=��a�rm(=�����#l�b,tuk�3)���!ө��x�B�s��5����X�	(�ڴ�E �Kv��`��I���(����-�����=�%z@sȥ�.9l�	g�	�y-<��WgԊ���|��������(����ÂA�8.W�W� D{�&@Lg�qeR�R�܉`pW�ՍH9�\�oSW�8�* +�޾��X}�U{�I�x�ݶG�h�,vd®s�vM��V��5F^X��T냂&z�Ն�7q�Ik��t��3
ISQ��Y:Uk���Y?ǒmHd��688f,wR�KE��a;z	ߙ	1-D��u
�!�X���X?f v��t�T�Y��+�`!�}+/�,ϖ��.������h����S���t���F׃#����׹��T	Nr��'��"�����#�@��v�UE��.�#3U$�.s �/׫n�?��-,�(�9��[�h��&��*��[xy�$���IRq�:��'�0�N�;^���<���u�A#�����L}�a��y�ܺlϔ���n�<�̢�ɮ3Sja��>�8�6�5��׮g%}M�G{ӓ����-J)�X`�C+�(��6s�Bj��a�.�}�QP~�8q_	�(lemG,����{��#�4g�W�]Q�<&*v��Yo���6�u|� ���V {�+��ǪR��k0#�c��*{��sg�ޞ?+�A<	IuǷZ��c�X�B��M��P6ݿ�6n�%���0�A�o����}Q�[��r��'^*�$&��1���^y�����f[|�5�KcUg��ݜl��ji�Zg�Z�U:`5a���+[��i�ciz��r��;����>y�W|'_��*B�`/�a	� �����yw�o�F�&r�G�gvR���(���c��@�/���V��.��X����\�-@+ܖ��K�]�+���2��y����f�	�#x�_j3�J)�Af�u���E���Kf�;gA@C�	9DW�¼5a2X���r+�<��;r�>2hW�ʧm�� �Y�7��4��m���L�KZ��S���,�,r�Pӎ#�X�s�]ˑ'�J���Yл�����@�3����7i��!@#��d�kPxW���Q�̟��u��������[�VZT^#1�I
�c(P%�6�g�my8���|$������>����I8].�i��47u�r[��pt��k�پ��j]V����(Ll�AY������08��u�TIT����(�{���(i-��m��n˷9��
πt���|����G����ۡ�|���r�q;����[n�.F+6_�_��%��O.�����B;���0Hږy!Ch�"}�d�Y��&֓[U^�U�����x�_���W܏K�
��V����4�?�xL�2%4�Yp"�T{{ ��݅�n��X�4���pr6>Hv乷�'��|57�24&i��;��V3���7�sr�.I�u\]x*J��h2�D�� Vj]������rK�\	��N֏�B5)�S��y��$E�N���f��uL�o5s���-����v��~^ )Anm��U�m��e�*��?|�8�$kOV[IQu�М�,��x�$S�]������#�+�3�_��QDzh���/�(ʎ|�c��>�L����3}��w����rPt.�������Ό8E�ט!u���?���[J[f1s�F<�	��Iy��R�O�`qL�)wy�Go!�~�P���>���t��2(���':S}b�65~�ÒcOuc���NM��u�@������J	��$HN�.0ekT$(�[����7V�'���^֋5�wʈ�@Q_	�}��LSFmqU��6�wj-�3Uܭ[�=��%�N_���Ej9ԫ?�~ɗ%�6ǅ%%X��O�g޳=�1�WG��4<)�s�	�`�znk�i����b��9'�ڲ���m��~�|�j}W�����O�OZ���{K��\����&+�{s樳A��Y��t��i��ց�+. ��m�^ ����1i����}:���.��3�4֡��7�"Eal^@���s��G���:�#p�/����"E���o&'ۙ����<;���C�g�B+}O����!j�s9��T����a�r%|�q3�)�#G��A8d��As�vLڀ~��1@�t͝�!��y0I�>��V5�~B"�j�O��{�w])3��oH����o�"V��j��̽����u�ߖ�R�MC5�4Z�-��%���-�d?�V��7����rGpL#϶\��ʕÖ�E߆s���/u�!�>N���Eh��ݟ�K{���m�o�>`����s�?:vЍ���[�VI����-�>H}jC��I[P�I������%DN]��i.2����f<c~�&)�s�U���dUt�֮��8T9���D���z����3�c[�0ͺ��iu���*��D�s�D�d�Y�i�
V'�9��FiΏT�·� o\`�0�|�����J���7fұ�I���� ��.0�d����a��P�����q�����a�E��)<�t���Ik%��]y0!�,�}O%#��P�� ��f���..�J��:�]R���� �@��j`u�aI4��%�c�]^c��u�8�GQV�Ƀ�ta�X�6��X/,mG�6�۷�Ja�/y���H�y�۽9n@&�#2�Tu���[�EO ��HO��;������,�5�������'b��p��Ǳ}f��"@)�W�_�tv��/��GU!=
p�o��o/�A[UF�F���eqx��0�3�;�%q$2��#M��q�u�� !�MS�z+YحޕKD��ͅ� 0��`�ý�kYDVѕ���L�}�RS)h#1}k�����/i����5�<V�n'��S����>�m�ӑl��T�� ��R-�����P��x���	n�S&��+KE���V�KU�!�A=q7��H����9v������d�I_�E�.cי���U�{9ɽ��Y���m�g�Y�������3?�T�v��ͩ��B��RexT��uW�N�!h��{$�j���H�4�m�I�_Y�m4�3n�c�������R0�hM�3�}��aP�ix�xSb\�L�G��J��/�čj
��%
u�d9Vh?���M����S�)�O��h<8?м^A��y�0ζ�1�ʤ?y�hn�����p��Gx���-ظ��9rCϖ�m������k3=��^ź�X�@#���)��w�'W�v�HW;=s�ǧ!���&"�3(�}F�NZ�� �~���������D��2���,#-��#�_� O��.�}�Q~�u�~).�-)�j$�OA���hMP�� �-�
,f��1d��#��ǆ���O\Ӌ0Q��vs4d����M���jsx ?��a��_�8�x�n�S���}���C;1��$�u����L1���5�C{�̲���;mJ׈*S&x9��T�;��ѫ�:��!RQ��*KV�]!1w��bO�W�%���/�>?�a��$�X~PՃ�� \*��3 �6;�8>��Y�'�j�Ü5�d��f]�	}���O�;��2����p�B��qy{�\����7E�l�/a��dFzi���&鷯�s��8W�~hG��GsUR���E�8�5��(�c�@l���}�0��-2�6�}n�� Q�8Ta�˰6/���v�D>	���f��;'�񟷺lU��J4]�����'SY<��^�җ��@�t�8h3���0������̅�M�ě1�k}�1^ro,2;����_���[ä�%��c6�c�,�d|�L��1�!,�ͺ��<� ��H&{�����]����7��3V�Y}���tLW�M��T���^�}E0�ʸ
z������!U�`�O�V�l̞�\�E�k<=/�Ӧ��s<U*�=O�tue
�ځd�������f��Q���
����%����{7^`8" i�d�.K�g�1��)u��6-7�޸eᖓ�S�:�+:���� ��;�����~ާ&�� sAQ%�K��D@�%��$��ƺYw�`(���������)��i�c�)he��6E,f��:���^u4'�D[Bcڷ�[�;����7w�%o�:PC}D�E�k���w��DQ���jsZS���_EKX��6g��S~b�SW4�+�	������]��|Z{nu�'�/^���fJ�41����cx��g��������O��m�*W<��3\T1�C�����P��?�YH��vm�_�1��m~.��P���^���,=X�M��TcD,�ش��Z���.O���;�Q=z����"�(b�~Q��f��FwE�����*#"!��"�r���~i��.���}���N�' ���y�iq[�#�~�H���T�e�R��O޻�&�����|�ŉ���p���&�]�Â �R��C��`��&�}hZ�Z�������g��z�ZJ��!����1Nq�K�O1�k���8�4ϭ�%-�"�y<���a5�?�$(C)O�f���F����$ x:��H���"p(@Z�0wS��?�l��Ha*gIa��}f�֩r� �ۉΎ��Zs0*�i�>E!o���j[�͹�,��\+6��|���r9�x�:�aڦ���XkІB����ӯ�_��D�^�nĖ��eyTsb�`$�d��刐��i^%4��r>[�FN%%ãqLNEi����u�X҂z����ۊ��Ca~TI_v��JL�Ү]�t�d~K)|dK���Q��@��ߺ�ze��h��u���
��Z��*����3[s��1˄��,Z�t;�?	X�S���L05�hb�R���ܟ_�Hv��Sv�\�F���t���Ki�F����֬�J|:�bVMv���#aj
�H�;��O8_�L3>u��i���Ky#�v�(�LXxb�n�g������7�7Y�~b�N�9%�w�E\��M�qs��p�~aUS�Y�_��oR�W�TX�	�������f�i�cwR�������1."���[��H��s����6�/��������wn��z��P�<�!�N���TA\�ߎj����[����r1�ty�{�"�J���Z>-*�h.=SYy1#���Y�>�L|���,i ['�"��z}ғ�>�gKt�2E
u���"�j�b*�v�<i%\N}�����v�;	mW�@���:���`�Z��B����m�A��3S`��G���'Up���r4�h�߅�!&bЪl�9E�J%+J���b��`���`�4������\+p�A�e�f#'�rF:F���8������rϼ�k�r_�+�JHuvRI���v/��=�Ua�R�ߌ����Y�Á]���-M�����!o8�Ɍ�,��&9h���2E����"�,��t*�s��]ܰ��{�8�aO�k����-:N������&]���4�ʣ�֐{�Ʃ464���b�\~u6[�{/�����D������k�׫�x�K>���h�-��ױsd����ݛ'�7 ��ע����Q�,��F+�vB&��#7(�X�"���	-��E�.Y�ƚ�G_}��t�;���F�4����uGCr�@l|~�|�.�S��K�&�\x�����n�h>���$R�5Ŵ����NR[w�kc�ղ7�j:)��v�fC-j7�^}�o9��I��
_g��?-@�m���2s9��7�}-����x5�K�4��B5��o/��,���.���9@L�����Ik�����!t�d�t��HŦ���h�]?&�Zw��"}��G�w5�o�kb��?؊�;Go���Bޤ~s��}�UYG:�Cx�e��<�;��F]��9�H�"�p���X�z�7nR�AA砽��A<>���r�33<�R��F��9�>;]�LN69ڙ�/��0w�r5�b\8΁�3DL������`?�r#"($b�����ʫ�I�kS�B��b�)nu���6+�+�p,v�Su�Ols7��H��=Sґ��ѳ?���ͻM�;�N�`����9����U@��}K�#�A�ĭ�1���t�E`�6m��E�~绦�i�ްҜ����B�>�ğ��P�u�p��T��b'�ڦI/^�\�*����=��=RFSt��-�/wV�6;9�P?c��Uy��wA������- �B �%�~yh'�E�[�����!p
����@i�����Y���$�K�7���.`1���I��T��G��x��R���J�&'��8�A���b����f~n�P73���d��c�H춶�m�~���Ӳ4�|_'X������K�+��>�}MV�7�&~��1�N�)��j5��C�\��D�wCg�8CYd��1�i�!�Ş)��}9�e@��X���Bń�N���Y�^�5C���cDh��V�X:�P>�n�i�&��W��X�Nf���|�P��00%���az�(�g�U�״et�*��S�yQ��k'�ɑǏ˷�!�ؐ�B�P��>���z�����'��4�I��SY�rB��c�x�
�7�u���x7V�Es[g�{�y���bZ6�7/�(w���C�<��[;�����B	���T������x�I�kp=��L��O�r�E�p<�n;��9����LPy%��yr"~��y���wl�l�B]z(�29��G���:����̢|*�n�X4	
�OB��>�?�#�
�R����ˁ��d��q�ǚ-�G�\A#�BD-;�Kw��@�FGRs#π�yC�B8�d�n2�?��TUj!�U�M�����=��]"�X��j�b�2���.)��Q���䫊.X��a1r%�Y��޷v�(<�6�k�Н*C��%S?���&�;
����]C3���H�#;�V!�h�@���|��Y5`�f5���"�ki8�h�iN&��dG��3�+I�E@Dp<T���-�Ć��(0������4$h�R��oۼv�u���s6�N�OsLskjX���!����p߱��3'y�J����-!�9{���9(��8���a��a�������|��H�P^�s�s�N钉��.�V���jD��D8�f��^��jmC4�i��*�"X���kM���Z�-�P{<�T%<t����
����ߐ
=��C�l�:<�9W�_6�b 
Q��["5Ặ��_m�*p��g�q�{��rO����wC�D�.8C2s�o��Q;�@��yq�*��5 ���İ��
hb4�xD��[L]K��+S}�W��A�.8����D�ҷ"J헵�:<+S)T�C��:�'���k)�ҙ�/t���O/������s��������?'�VCUul��c:V����t��_F��R
��b0�ڹ�u5�F%�b@���C��>��)�?/�ET�z����&c���29��g�߰�GP�4y ���
�[{��En�َ|}TJ>X��}�xZRIPaxX�N��J�*`v��˦����bvZb�A2TN.�v�E)�ro�c���u�m�)�	X���u\�ؽ��k�7�����<\`�Ga]��P�f)�.5�~�ލ��΀:����O#J�"��gl�^��EP ����"/Б\|͇���Yyvzsj�r� ��m�8k��d���M�L��x�t(�1��-O�U��!ڍ�Ka)�^�;2��s�1�yu�JCQ�s2�ɍ�%)�Ё	��O
D�ϔP�J�j���m���/����k�.?sJ����NfʸX�3�U�����?;���X=�Fn{�/ $�	;��v臧X��ʶ�Th�'Y�]gn,�f��.��39�G����D7O~Y�T�%x7Z_��-��20��~�~�YH����{'!�m�m5}*���oqV@u����sA�2N��sɱ������q������?V��U�E�(4�(^m��䨭�?3�l�ntc��Z��{]�r\m������������g��J$TU1<C}�A�@>����L&�ǥ�}aa��#˝��~�D'��%9���c�W����QS=�I�JE3�R�+ToM5x�=l�皡��:��4�����:$#���I$K��ǑuM��@���#o�py�I�u10^���۫�n��ֈ��!�$##�v�����c����NN��k����*�b��3_��P�Ζii^���3%[�4-����0A���f�OW��AX��C���f���~z�e����K���F<�ݺ@�ɡ�&��+q�&�|�wg�g�]����$�eyv�`�Rp���D�Tq�k���|N�	�(_"���&�W7Y�Q���dY�Z�R"ժ�G�q�>qӝ��l��j*��kN�:��M�p[�b��}��5&/H"�%h������s��U�ܦ��r]��v��J%܇�a���kB닫�Db��j+v��G�y��紿�NwY�OHu�'U����`�Y����F2���@��$Y68<�B��*v�?�������g�,���EӍ�&!6E_z$�G�}�����Iފ�&���iw��������M��ct#ҌBX齋o5��f����Z'��zQoe�NP����+��æ�CaQ��������as��[��}#}���AnU@=�$)��qe����,�?�fR���������9�o�8k/A��E�5��_9R��s[���\$��_D�s`���(Q�a����,�T>	<m��fp�@��}Q5-d�#N*�6.�ǃ����N�]�2?q�R�xI�^q�b���^o�n�{�Ϳ�<6�J�
�(��P�	\W�bU���f�j�9Vg��VOç�>�t���F���{w8s`��͓m�Mb{��2̩�q�4X��'2*R����U$r�\*[@ ��gCux�[�`����E,��0G%k�q�j�Ԕ%���*`� ��������Z~�	F�@2)>�-
6�;5��djfW���6��k�@���討�h��˒#X؀�D��S���5UR~�6o�i��ub�Qwr�zK�{��&���2�����wq�jR�BO����)�-O$Ј�h�ع,͇�ӓ6y��s:Y����@��8�����R��=*]��T`� �i�օW�2���ih�MBE�I'$e�E������p�H� 7�G�f���>m��j?��.�\ovw��L�����=�h������o�`V���~��T7��Y)�y�1�t��q�u���r�Ɨ	��Ho�!�VI��A��	v�o�(�'�UOC�σR>�^_�����ivY#�|�[��1����?�g�mi�z��b�,ĪaeD〇o�9�B. 42�4����(�y�UI��}�n�ԍ60���f��W7��b��5��\'�0�/���x�i�G�ۊTksC/D�,�}hq�?�V�<ƍjeN�p��SP଒�m���2�I�D,vR��eԂV�����ö^n&�5�p.�:`��S�R4m_��H�Ѵc��V�K���w��77�B��L���9,ړ��{i�J��0��o+C���~��5�H����W(�I�;>/�^�N&�)e�6�3�B��`;r��)e3��)$_���R$bX��z�w[�+R��6��s�-qe���*G�����6;7�.��N���J��ɒ�XJ�Do]"�O������u%��\����x�x�׃�;�JP��?���n%x*��7]Z��@���XS8Q���c�az����f�LQ�ե"}}\"�^fo��GN�iaa����}J�J�x����x�[F���	�W_���I�Zo�z���H4MKj?�E�iY���q�M+�k��7h������+ݴ���hA� ���FX�l����g�!�2�$�j��!-��`��D���T����"��ǚV�Q�ܓ��2M���Ʋ����\Pˏ��D7��R���e�Ҿ���/�+��$�d6u����X5FK���[��h����Q�Nn��J���]H$n/k���v�������>�t�cU�#��@U;������W|�V:���U+?D�&w�l��q���fԩVl�NF�Mdf�ռl�b��i4�Y F8���,I;��[yT�~1Y�����v��r�����F�����䴌���Fu�$�T���[�m�e�����[K�_���Y��`;^��q���������n�%Uo�9�o�z����VeFbw �x*�r�O�n�!�y�u�-�L�C�:�W9�����ʊC�H��߼@'����|k��;�tb,��fb9���:n��F�"m~"��]��������(�*����|�G��ms=�����P�$p���T�:�e�\�_� �ݪ��M��▰8%����z��l�K>���jc���^D�_u��T�
�3�>�\�3޻���^�j��N߬�X����!
6�^lظ�uN���e�r��P/�����ڱ�_�gbP$�Sx�Wg.,�"�����J�
�Ϯ֦=`�
kc$Ԑ��w�+�����
k��K��Q�%��nc5�!.X�M�U(�Ѽ��+�Ā�����ֈ����� wM�[���
n�a>Ɣ6&_C�D���:��?����6N�2H,��J���� ��i��!3[������b98�����������C/���P���z��~E�9.e��Q���Y�(Cwvɭ�̎�r���x�$�p��a��jX�9u�N�=bH^ �����)ҊR���B�,vl��[������;����ϙ!e�{�ɖ���[/D��K����k\g�%#*��w�?e�#�p�����U�:(��k����l/���#���/�Z=&���8-WB��1���x:9'D^��rYưt�V��Wu�[�ro��_c����d�����/����R�گsO(0���#�7E�͸69tN��7u���q��R�v�j �s~j8�	4��� J�rP� �"���d8e��]d�@��jSq˄���F�_����nTx����ܳJKh<��&��2Hu�J�3:�#����HO�oM��,��R��`Π?��(PJt,?����fnbLb��H�����<�`���
�
(���ȗD�[p����u�6��������s� �zV�65�;jd9�oM,Mg��ɥ�����s�v�A�c̯���������; �}�Z�ǫ��|rd���e��6��Z����xQ(��<���T��)�)���HOq����Aqe.�ߒS�Gfv����RXJ
:1���\ߏǵ��(ʸU���6	�����%�Ct����8q�sxB�2"[~����EK4�z��=�f�������ʎ�)T�p�1ُ�� ���1�CY*rp�a�cu�������.���EY��BX��7ڍ��ҭw��i�(p㱸���S�\��+Rt�]�-;�kH`��a��%E���=/T�t�����/y>���9�������rm� $��_-o�:uF�������Uw�A��I�>0�������=��M��m���ŀ,)rP�9���Ӹ��2~����=���;��[WK�Mu���*^¬�D�#�p��JኑE�����N ��yL���|(���V,UB���Cj i�<8.*rg�0�m��'��|G���=}���h~��<a�l]@k��:���'�7��R���b��h�A"�#_ʭ���_gnҪ<�U�tVjى{XV�V���w����o,����G���{�ϒmz+�9�ƣc�كy����wO!�mz��+W���_�X3@qV��s[=�H8z0��5��(X,�L@S��"�X�}H ~�t,�D�d�kNmAu���q�)Ӻ�j�,±.������bΠ��y�u�"��-830hOm�|T�	 ��vDۍ @k�'�m��ǦM��à�q����������bJ��l��[�$����r~��H1���˶d!��`lPm	�]�ut����o�Dg@��}<.����9R^�y��pM%W�Y��b��-���	H��qF("�Z"�-�	v�H�zt��Y�V���&ó@Z�I��{�j�O.���1WS�,.D�? {��HԆ������׍��?oH� Q���`���y��������0xN��KE!�6ҝ�Z_����j��@�ذ��U����ZWjGC����f�X�d����Vo"Y�xr��C��^���ﲣ��&e�YCJ�@���:t��{�7�ԏj8�S����GUM�tf:�l��Z����k�S����l��-3����,q�!��@�ɱ_k��a]J�Z«H���1�rpJ��ģ���e%8�2e_xD���o���������W��b����_ݫ�Ti�������u���S��`��*��(���7��ZW�EtD�à��4�?9ܧ*��}�ΐ�/ٹ ��N~ҷ�-pG�#�{�W���������+׵�zL���1J�4s�q�ի:�牥���Zb��Ԍd���!���')V0�s�(�`J�ņ�<�NPt�������iVX�����}�k䶓FV���3[nz��޿���m�9�5W��0�s������Ɓ L)�èazӨO7.~�U΍���\&%�=��9�S2֨>��>z��l:�/ԫ�zvQ�π��`L�>����[�ͨs���dt_6�u�r !��=삯Z��ouuSA�=hYo�<��a�q���+��H�S�I�Ɂռm��4ȥ+cro�����|�p��>H��'ww�I"ki�����~���Բt�EU��ϒBޙ���9%π2^���u��u�PH" ���=�!$)�-�E]�5^>����OP��������X��֖����"�uQ惍2��/� ��XE�n�p����{���(�t*�m��R�����������e$�T�,�����"Wҵ�B�H���|�98DG$j�}?\�x֗W��X �����&��h��g�@3ͤd��D��� 9KV�;�0��#&/,A���p����ٳ��DЖ�'E��4-����}Ň�("ZVs����Bd1^���.��]�˗	M`�Sx�רU�m���j�l=�Ont���S���6�"E�#�ĭO�@�_b7�����i���`U&�R�����@�?�M���a�������p�j(�	Ә�e���gou2_��}{��2+��B�C JՊ��+*��9�s/� �����0QUp 6m�Z��
Uz+ ��M¯��ڶ�3aLIWN+\L�kqȼ��P������R�M\�'��[�U5�����m'�t��w�,A�Nq�����\YUB�2�?�#��}!U-�YK����b&�]8�n9&A3~^e�!l���rs��mx ����U��yug�)�g�M�e�2J@�0g�^X"��gЬ���?J����~-�w�>Շ5A�·�Am�	���Z���W���ؙ�]��z}Ap�g�{6����`�蹹e���B�ǅͧZ�s F��oD �6�bH���ݍ��;1�@j�bE�����,��){*:���}�As�X��]]��� @s�05�x�TH��%�Oe4𩢼�5Ģ�b���I��wD�N޲��O;(~qcYl}	$T6}�-��0���tωv�����_����Ua߀�^���u�!���8C�.����� '���Lʆhz�;�v�$�jF��G ��\C�<	O�� �:��K;m2
#rȘ+n[����z|)(%L��n�|/(A">rB����C�wYۗQ��UM�j\O�lq���fݐӝ�������<*6/�����Þ]'{����%@z#_;�ڱq�DgI��G�^�𕜔UX)�j��� ���E��{��ԛ�L��"�t����ȝ�E'B�}��_��V�%f�7�k����xl+�b��'�!�<�ɘ�̶%���o+�!X{|?�}�.$�552�C_U��B-���ct[s�J���{�N;ۘ%&ro�9;����sk���S�w�\����IOMD��R�)�`���((}GB�i�y�P��)�/9�����r��k?�t���r������kG~��)$"�q@���Z}���ei��{�0ߖ�B*�%�mG�Ȧ�YAN����A�*��� �4��?7��	����hC�ýmrj��C�{lZ~h���A@���\�$��R
`�$Ϩ�ufJ���>F�ilx�H�ou[�(��p��~޳ȴ탈�d��;t�l�F��"��5�h�T-�E~����I&�C�x��ɭj�_N�����>�|�j��wx�/�[�rۑ��>K[g�ްET���R��*�����&s:n`�Hw["p���C$��
R��2��9�K��5:W�HA5Lb�B�����dۮiI��)	1�G���P����_y�d���e)���)Z(cX����x��]�+*��(݀�4�z]����{%Z�,-��"FFG]�Zi�B���K_�"J߸ �
@١������Q�甮�mb��үxX-c�g&��W��kۚD(�%[�X���"u_4�����h�̰@�)�D��Gp�Z�Q�4e=�ؽ.�U��C{ҽ�=���Ӳ��Y[�V�q�2'��zF�31j�AÄ�4�>Ī�pV;���`������-�����U����w*�>�'W�,e���M&j�Q72�Jc��d�X8�!8�S�����u�����1`��	6Z����8�|���
�Jx,�=�,'�48�^�� m�A'��&8d��FZ��c]r*w�z	�R��n�<\Љ�J��ݙ�xٛ��x�*=���H�rҊ	KF��	�Ru*s� ���T��1�5��	�t��9�:ᜇ��?Yz�U;���[;r�7�Y��[n��U�K#�-b�?n����
��m���
?�&S�3�"J$c����NMu�5Mq_J��!9=�\���1^^��h�����9�sF��z�ex�|N���?�L��!�����\��K�X���r_��]a�R�&bB4O2��G�v�v�`t1�[<���,����~��'�N��B�C:�%^����A�C,��c���T���x	fֆ�MA��:�.�ѡA%���X��XEuX����b���e��ٚ�HML�Vc�F�E�:+6ss2g��1�FvH����N�M�ی�#d:�ǯP���L`M�j�.����=T���\�I�W]�IJxW��Lct�^�O��Grq�ŵ����<�s��x�;�hEM_�7���}�DX�f�D��]�͹O_�L9���-�둬e�����υ�fNV�����Gu�J��Tm�ث1c<"G�,sD���n����Пb��_��3��8��D�8E92��J"O������I���yKdGc'LT� ��Ҿ�0t1����k���I&��;�`!OX�7��~�p��_J��RYl[���������k�J�i��͟�ڐ�K��'�~�O^�#?��OmTu�ww�TW�߯A�d㣤��4 ���2��7���fF=B�����,Ϩ�-�䝂L���M�Q�Yx�#�H�8D�R����,�i��$�̨�%���zu�'fi 1�G?���!)�Ք%^P�r���"ӂ���x���P���[�S��Y�*���~�� "aH�ɑ�ڪՙ?�(�-ړ9�$�ȩ����8�3\�Ŧ	37��U(n$��O7�B����^��q��.C�|h��h_���{dJ���Yv`�$x&0P�V��a��D����G�6뵕«�+ڬ�@#��Gί�ѽ(��y�d��yĦ�>��'2�51�y'Ļ]=YF�a�..I>���Y�'�ǖ��iz��	�.M��4w�D�-$|�6J�}�Bg���(�:����j�Ԓ��dN׮��|�f>�zZ�K��:I
�b&D�g�i� �!���k�S�vFJ<��Mc��R_W�,�n�2���$ ���Vi��*���NکKi
8E�߫��#W�a�i�e����F�v�`�u�Y��F�]�fv\8E�����n�� ���!F�gM8���%�b����;��
���4�i�%"	��������M�N3x@��+�~7OȈ'ۤ��2��~ݬ�)�Ze_�Щ�{6�r���y*U�n���¼}Y\$��D��"	������ų �û;U�C���f���%50�s�ДgN��r9����L�!�-������?ܝj@;t��H�-��*���|�#�||3!(�뿖��G*ɀ�E��Uk������s�u9�X/�Dp�z�%F"���`�]hHqE�j�U��q+��Zlo��/J����;d{�Qi����R+�Z�!f5�v��=��;�ޭq��c�VB�w�ITW��.
X3�=���h�啎Ϭ�K��-���O�L���͘׆Xx�dQ��a6s�Bm�A#�VL��dyCb���s�ld��Wr>�I)��q]>!"%{/���¯�?�)Ci�9�F��pʬ0�gI�p%u��*��χ�I���5?�$����t�m�yC���pF� ��X5��ݗ^閗dEE��{�Lj$�iʃ��n>벅���u9110�	Y=�� �6��s;��9np��I��� �Sӷ���Ua��&�f �nhƖ֪����v{��(��3�U
�s��y| �o�����ۂe���%H�3H�����2"�4r��g��RX�^y������c||�[�E�j�(U��}|��������Iݺ	�E���;q�Ƃ�vVZ��[��c����E����� ��~Sg�2�G���D���#%�X4���R��Q�,�m�շ���^|��4�Dyf��vV�Uxٳw����@����,�����-�
�6E�7���'�<xb7������R	���摶Vcx`,p��	�߆.2, ���յ�{�I@�Z�.@�܇��.��������O�4�q�A>py���j��J_R�%��5��&��: �V�
�����BN�����C��~(I-9*�Qk�/�b�3zU�-�DĐc�P���p��fu�^p�w!�2@8��eB�nl�#&tA"��}�+;\N��!�Ȥu*��t��y�.��m0��l�j�KJ�_`�(�6����0���	�@rE����	��=I�O��O�������	1�s��>���\^�\�f�T5tU���G�?�t�	�w`	�t�'J�Fj��n#�z(O��5�$@�}XHtB�k�;$LA5k*r��T�3왪�D��������鋡Y7��&�Gu(������6�%���
�2���/O�:l�+�.YX�s����~O2�˲Lz�hQ ���:��0���:�[��G	��f:�'�Bu'%)%���ɓh~����Iu}�rJH��HTP�������J�p�����`�
�_�*N���F:m���`jɛ���b���U��'BZ@>DCQ	���_~4�'ޞ�G��@CN>���ʄ�:`��Cd���$�����
�H�9J��Ʊ򂾋�]�����J:��Q�J"E�`���-�lw��B�-��E�Κ`¬jE�o&�zMx�Rb~6���6^��xe@V/;N=E7��=_ہ1<�0̘�EՆ40!�⹨8��� 8�؃�اdd��7��<�%h���٦p�u)�'�+���Ǻѭ]�cS�AB��kI�sȥ����NF^:Zǖ�t9 KQd�7���*�9N`jw�BQN:n�-!��m@T� �f%�Q�_Y�e�,�W�Lڿd�t��7��d��r ��S�3rJK�� �rӢkV�~����g�pe�7�"�9�>=Hx��8<i/��CZ�Ǝ��(����Mm��Y��U�7B�Q-Ӛ禊0��n����krXR��~�L��ƥy�o�n��b��zC��f-&����캱mO?a�k\0~12���Xo7�1��H�W�9*�*+�>l;0�?Ju��Fl�[$��9��K�j"�U`5U�*mgoȪ�6��Oҁ����ĜpQ-W	/����}$|z�W���G��JRr���Y��4p�������&���b��eo��M������&�B¡� �P�ę2OT�:g�"�8��	���/9�N�N��R^b�e���L�!��r ����l��t�۽R%�÷�����įHx�_vg5/�lߟԣoaό�kRC�bFi����z�0x�0��
�:��s��� �۷���w�*��rS�e@r� ��h��C�V�tGw������|?�rI�0��:��
ÎS,Q}(��aN$��O�� ���DL,)��ns>}%ux�`zQ�I�϶T�����1��G�Mu�e~cp@��9�{<ה��j��s1��(�+�v(lYE� eg������R��]OZ��`�VG��0RX�I�C܄�p.\@%�`��n�{��>�9�Җ��)ߙY��X�P�BM����[����F�W+{2��kl��)��+��}úw+9��l��QjIX4\�Ů[[���i�â�l��K�<�*Ps���Q-%^�$Y�\0������#�����L��!k��9ߺ��K�
^�,K����QVਇ	��N4���R6M����>JP;�&����2*��&8A��	(ls�E�G%&�}^��OW��yV˦Q�OG�@U�O)L&-��?�)���q�={'���R4� �xc�%m_9�����ȓ|��b�I��K����p�X�:p�3|㽭;@v̀����+�j�+�B/~�~�;z���Ikk��UA�^HѠ	�a5��E�Ư�F Bd�c�`Hg*K�V�R=6���̚��,c�����>�<P�Kq����xe��@�����RZX��H��"!��y%g)����'���zJ3A��=�H��m���%N�-�H��	��KjO���߁=��ώ�X������=/wWz,�|*��0�ň95ݹ[��]z���)�
?cm�R�\
�Dv�Ԏ���4ċ����iU�G�ʲ���>�R�y���#	�����3� �"�0pa���,�Auy���a��o�����u6��Ѭ�7|L��h^�QeB����S{�:���sJ������odz��%9ޔ��ԍ��IST#b�����/��]ʜ��B4���Y	��r !X�@`��N�X*@� 0�F�˴*!"r�Ʈ�vHv�#����{[�YT�a1uM�0��8���T����d�M=�ʷ��Ը"�����@2���ok��H���g:,�K��؀Z� 	�姖<1Dz-Zz�o$�����T���$��ժ����U���뤻	�Sk2�o���ZC^�~15=�����G*���su��-r�`�,��j�E��ܻ�B���M�I%|:�ފ��f=m�gN2��!���{m��4nZR�����3�U�ҋ���0��?K�����6�KV�.�>��/�����A� >��b���X�60J�tzO.�7#���"Y=dq��c��.|�Cz��k$���t'I���g���[nh��{8�?��̏�CDb+�߳����#i�;������{n؎����dN�\.1X_��t�	�
�O ������!!��
�yq�!}�!��Y+N�I��kS��?S啝@����h� e��J��L8�:�lb�S��5�6���ML1���(H������n�vWX�1֓�|!��J�$n,|�_� !w�}�{�7nif�4^:1���'@�#��Y	�5������ZXN��`謔H�o^�)��&̣��|oS��s�
XM��[���;KH� �I����<K���tv�H�t
5❓�`�-}@΀��<��ql.�῕�	���Qj���ɼ�x��?N���&l����B]��p����.3*y�4Z�����Ѻ�ƹy�K�K1Z��!}T�;{��� �9/.��
ND9�y�v~X�KLl(�t�&ح�MZ:�.�y)^8�
?Z���]t1��>����M����5���x�y�x2֠�a*�PM��:�D�z?� Ne���Ѓ�x���{<��x�|'��%�Q��Xr%�~Sh�Ta�]��R57s-�88���q)����b��c�x*��Ӎ����N�6���Wש�Z�G�ꎥ/1�5&��f<$p����~� �HV-<V�M�q�X���C�)/��0�3#a����e�<�r�7Ź~
J߫�6�j�� =�۟�q�È����R}a�"Q��!ɚ�r��Z"La
�Q���&i%�[Ui�.I 8LH_���z��`�RJ����=n��� �J��p�f,>����A���L�פ�|H�'M�V����!�|����������ϴ��Y[�/���6�"��	�Ոr���CPG�$�+�n��t�
����RʞrW%�pY�ה�uQ=g�h�"%KJ�0��|��TbC�	�e��n�%��z�ls����N����f�m��@A%Ǒ���Hp���ӱܖM�8+~&�@&��⿾��;5�7L����,l�<G���P�Jw�p�y�on�I`���/��~��ü����X;�S�$�Es�n�0�	���Y�lG"�wM3K�Nn[�6!,��~	�$Ub��ZVNuJϕ�,�8yY�'��ⱏ(K��� B�Na�PҬ�ފwpB�7r!�$�`0�t�]�6��-��y�tm]��Q���R4?q�����R�W����.�d͂xE���?xk`��O;YM��^�,9�]�M>���X_8qS�~��),�s�ޒ�!e�ͅ}D�k�Ƃ���KT+�
�Q߈��h��'�@/�e��XU;nx�a021f	���~�M�wX���Z�Ql ��y��5|��OCJZ�&��V��!u]��os#�_���c�1�v�6�{ �����4�m�X��Q㲸<� �(h����_D&j�9�<���U���f�@�<��R�0#�qrEb�+���?�}�H��Q�{/����֝1�[w���)�����NiC^Q.L7R�,/�Q	%�Z��\ �x���-WɄ-V�|��K������#KL�����u�qa|r,�p�SRDPhm�ܮ�WCUur���f( 	!�h"���7���N
$wa����v�Z�-���;I����֬'�nE�����1���$�8x�9�����s���m�����E���ѓ���ؤ��T'���[��Y��7W<v��°��6B��:J=�������(d3��Z�䐱um��
P:]��jj�zf��3�!��[v��@��D�z�'x���b��D��3�'��|	�b��Ò����种2��S��\*TR|�P���7�4 �e�����a���z��7�?Pw�ƆdN�<?��Aŷ���A�K-g�A�(�Ψ ��|�k�
/d���?y���� �B���̉r��!��s�d�!f���_<E�V��KU��ms�󽠕EZ���,���yܠ������_Pu�V��j��dc9�ҥ� D�Lț�cl��.H�0�%G���{q�̦l�`�+�Z{8B&���4���L��q�]i���${xY'.6o�)��-�n�B��ĔfY��GA�Q�O�`�v���ig�V��ܮE�ak����0��a��ս�)(QR���j�:+�%,�#�ʼ���&��Ͳ�>MV�4�>|+���}�.f�؊�l�]�g����o(B�>����W&�jh��D&�ȉS.�#峺$ӢI:�*{N3�?�3��cA�����y(J��V�6,�@ظ��V��]�ڵ�����p���Y6	-yl�'X�X٤����h��X4▞
3�d�|�|��1Ӭ�]�N0����Q؆�4�W�P� ��c^��g�( ���щkC$=/�h}�V���L6�!�I	;+�2�̮��
�-AE��Ɠ~���S�`ӳ��G
�f5st
?��;r�x����F,vA����l��#j����2Er��5y�y���j��# d]a���Y�"�^����`��U�zK�%i���^�,�������}�ʣp���}Q�t�8r�(�L��E�}����Zb7NO2�����F	�v�Wk6.��05 �d��P�p��j�ؙ�!��n��xڦ�����5��.ͦ�#����*���`�Q�$7��䮁�mi$�W��`�����w��s�6�k�ia.EtECx��StɁ+˄|AL Ȏ���<�=���eմC(��tIU���䜟W8�'�c�U27 ���`�ź��,!K��İ7k G�O��� ������@����0����(_z\�(�6���r(cX����6�q�8���5�3o	�(��\t�k�ے�֨���o�v�l*�`֔�J���챎Q���a��y��:���>�:n[��s獗;�pd�0nU��:%�.s�U�6I�cc�S��5�
Mq�p��A���(iҿl�0|�>����L�sW#
({&=���jƚ�\�M�j'f��B�]���URY�
^�Z^y�PǼ�K@u�\��D'9p�;�&����SJ���,* ��
q���8��m���wwwd�?L<_r��7a8X�,�*r�-�T����Y��R�y����t<���빵" t��� i1�mFt���9&��	S��B꠿�X8���Z�b�r��U�:%�/�Ҡ�L����=cD�T��7f�ڌr����yL��l`�d��E&t߆���kY�[S*Y^n�Y�6��lm�814�59��7��}�ޙȅ�c��R�uEw��NC�y����:�^����@��L&�9�s&^��ݹ)p���8)�_Y�Qc��=v�$1܆���+�鮁1'Ht��j��|�0q ��.����a1���T���1r�L��� 8��h.�ٕ�Y��[��X0Y�Ë����_E�T�1�,�����I��FP&m&�Б:ˈ_v��A��vc��
N��(OQ�Ў>�ێС�?U5����3q育��Iؙ�dnN!e�\3[ɟybt�5 l�󊥽�'aZU�I��:���$�˙x�[��Ov�B�a���G���m��5�N�F�e Q�P�ǽ7�%}�:���2����&Oa�x:�wq��[�(�˷ՃCI�ǎ$�T�?+X�y�ՠ����	����d��!�P.��Po��%���#w�o�L7[&mrĢ�;���X���e|Y�Ti�R(�Y8#j2ErX�{�?Rh�	*	�fT���#˃�8첊����7�����˵�iO~�v��3u�k��ç=�����A�d��F0Y�b��{�q��p��  :�![䙞J�^գ��L�T��۝���$ӝ�'~U�<�|OD�l\l��Y��ތ-1�q�~��2�V�T;,A���\z�;�\\@��U�hÓ�"��Y��j�״�k�K�z�ݴ_��YAGL XB��4�l��؞����~��s&��t�(������Km�.س)>�%r����KO�_���%�]3����:��)��{ZZ�����xW�K��$*��e!;�)$eo�!�+"iIL���#��<}�/z���JWCu$���\�_���1���o=&#5œ|�"!'}��̞���@��?�b,�Z�aN"��6����V�ݑ�y�=[[��
��3�mX�Tc	\�>�8�s����$ @�:8(G�y�r
���ZD��e�Pp���d��Y�a�RI�'���3ib)tb��]L�L�ﺓ"�2��8?����O�������3Y�,�H���
c����%������g@������� {m�Q�J��%;N���j�<U�����e���B~���&�T���:2�k_=�.�f\��*�M� ��ގ(<�&�~(�	/n(��ߘ&���M��g�!����{C1����
HF ���1z�����Cf�ɵ>y'�U&��-�:��n�bE ^��V���ݒ��W���j)���4���3�]|$Q�4C���7���G�DӐ�)+��ԏ�O���֊�ar��$��2U��������l�;�k�{6�^ϝټ�����5H��������!A��A#��6�`�K;��\Dj#��K8�>���}�'g ~U�����Gi�c�u�p>��b/b�� [n`=Z >^~�z�1����ӭ�� �}���BL�CoWL�cx�̳�}�`啌K��O~�i��ŷ;7i[��k>+d�7���w������O��;�TVx	:���WP�%ik��׻��y5??DP�p����͹rU%5�} 3Ra7����&u����}�6M2+�᪇�q��o�3M��n��ᘬ
�X<�J�*�@�P�+�Ⱥͻ]t�x�o�jWG��q��p}9�]��
��{�=�m��P�Q�G��<8[K��V�Q����ƻq���>?����9	��c��}H�n��f�\�tT��Ja�a�B00�%�ֽ��D��_[I����r#B)&w��$@1J#gt�=P��x��˙���Ӛ�wpz��������}E�/�����σ�3����m1��y�K��O&(v�i�Z��P��$D�H�v�C ����_ԡ= ">���ΞHtZ&���w���GR!�X�p���9��ao\C��{Ѱ�=�_e�R\hf�o��|.�fUT%7j��"�6����+gv$�Br)|�:,�S�Iu��gC���"=�Y�:��6]�+I7�-��k�,�K��
�h��v� Z����qӊ��Y��r��;�m��Mt����Cv��E��09[����+�7��[�W^XA;��)��լ)�3H�/9�X��7��D�Y6�,�yO�}�B��/�*�\k���t��l�z		&?�3A�7D��=�^ݪ;������?�O��y��l$��lo�5��K�;-饻��N-F{��Yx�3���$q'�BŻ���E`o���s��Q��V���װJ�C��+04��1� �=���Zj�6S����a��ӏ��ۑJ{	?��<���J��՗�gu0���h�H�qC��2���>�\����ꉜ���X�NnY����JӚl�Fg��vNMh��Ly�ch0޻2?V��� � �U�\� �^�TN>R�)�+U�}���fP���5
\	3�6��<ʮ�Q��`�/�G����x��b(���'.��2y���4�^E~*��E�`lO�,�-ZA5傂
��-�ʩb��˳�kp�-����'�#m ��4�&Ņ=����ۋ\	�Gk� H�G���d4s/�ּ@vEDؿ�i������
p�u��Ӻ����SL����U��F�X�]72��9�)�a[N�'��+G`��o886��S)�g�z\�%*)��~�ĬU����v��3���#:tm=7�!Q��Y�	��xo��ՃX ��[�2� !�NE�J+������IX��ݯd쁽"5>H�dW�"�����N���A���kL�.����;	�i'(K# P�7�g��|�\��3����/YIWQ*���:�t~6���i�g��>�bZ�=Pi�/`K�Z�Q�E�� Q;}�B�m�Y�sUq��R�J��ڲ>�E�X��d�D���I�?�{�o���n=cSf����D�l��tg*�b�n��e�),R݊5Ą��É��nd1��!$r�*�%��r��4�\W���5a�n.��)����(�z��<�O.5�m;�{�@Z�7�GV>1�.`%hP>��`n��A�k>3ň�#a�b��x�>4�&z��b)��������%1A^l�(����ү����������4���DJ���{�ap�6����\��k�o�(]q¾oW��Qx�_�E�h��"�1�k)��4��c8��H췒�lC�<�_����I��H�z���w���O}��<�l�&|� n_�a�R�|�sd6. O�I�̦5:r�U� >?���)��~!�CZ�Ti��}Q e�)ַ�mq�Y`����v���˳��"�@��/_ê��x�-���zD���8w�>�Z�\п�c��ɬ{U��U@u�k_�j�-��37)�j����ʃ�f���)#��n�jġ2��]��|�,#5b�D�Q 0b?9�Q�7'�PXU�k��/�^&1�+�{��[[T�D�p��|��µ9Ƿ���8�,Q F�i
�ElMW�<yU�+���ޞ�5+���Xi��!��΍mo�Y��-��x�uQW/�y�xz�u(�K֭����oDT.U�Qi;[�n��ʑZu%O�\��v�%�e��A4np��BQ�k��?�_v=�� x����bشZ��V^ss���YS�I��NE8�@�{�qg���A�2�l}�R	B++�iK^^��� �j��0��~���y(�~g�7���ݠ���L�s���Ih�䜩�����9� ��l���o�J;jM��TmExSk��%����˂����U�dh��0�,pM����r[�:���KX�`�ԁ��Ĳy5�x�<`�oץ�͒Y�V��k*Blh��:Jx]W�|��#fl<�sl<�'秲��~q\�
����N�lrr4_)/w}��7%��A;<�e�J�]٥�m��ob���9��⍃��P ��<��˂k���N:L�Y�eH̅[l�x����:����I,M�De�?W�8�5�#/�ND�Z�=�9�N�q�^��jb��&���=?��=4WO6ǄZ$�\Im!]�[$F��]uW+#jƟ�Z��O�).b�����sd�,��꽻��@JE#T�V&���B5R�SѶ�Ӓ�|k��Jg�B��q^7�K��8^�H�3�A����X �\�/���X�Yy�� 7���u�X@��V(702"8Mn@/�BS�!yz&S�M�
]��̇0��Q1�~k$�֟�P#����,:������H�V�F
E>4���i���(И�X��eg�\�b,�:��:
���Z��ۻ��������XR5|�s���q��	c�A�p�E�g��Q�����Ƙӽ:���I�ßi_kэ��#f�zV�g��_�{=�^�se�i�\��y���~.���7����~������7
�;��W�����!R@ ���jbl�@�:�7�\�5���'��γ� ��7}8�� ʱi�Ą���&\��M[e#s���Y-����f!�=Դ�E�K�Mi������3�T���e��s�ˢ�H���@��i��~�WǠn��բؓ�V�d��H4�QpƎ���?�hy�������!��������P�ʩ[!�"V�;ԗET����*�
��
�W&`E �θso��7P�%aO��w.:���y��
� �ϊ����ժ ��N�<�\�)@6�]b9�u@���:���,� !�,y@u��d����r�ٲ>:R��ЉQ��g�2��׼��m�c�	�� #����%�e|�\�<��Ä�&m�/?��9�,�ΦmQ4Ơ�ͱ��z�T�����]gq�$t9k8��LjT(����p^Z����� L̫`�(���9LE Vc���y�u»(#�ρ\Q�n<1Ǡ��X��{���a�S� x�dV���ɘ����0w�}'���Y"�4=m����	ø���6��;?O�14:�!tb��\Vv6�P ����t�z"�!NsҠ��|Wz��S�N�eJgOmP.���ixܐ��z���mˍo���p�d�`�8ӟ>^���,�D�J�S(Lpj@<#o��xfj
{���σ��׵�d��?���2kSŕ�[�ÒЗ*�W����}��>�O_G��$���[�A��Bu��+Jp�Ɖ��x�S��e��{��.4��/���"��H0��׺h,�)��ɿna�r���1���j�x7�6�J�dV�ktt��Cǚ�{6/��㾘_4M�A)��ᅪ�ߢ] �h�����9N2�|{���%��=eU@ɛ���E���Ǽb`p\gj�!qwˡ�jx�?���՛��bw�]W��N��#�-��X�5{����v� ��4O��*��Ow�?d���XV���]�J�Ȝ`*g�X����l�=_�H�HA�mi���3�lC��E_��p�Xޡ!i�f�P�hg�l�(����mJ�B_����~^��V�5|ȸ��]EP��;�z�q.v{�R�E^,���{K��2BT۸p8q�t��8��S|x/�g[���3��1���9S�ɜ�fP̘d�Sn��v���y��ic����g+f���&C�:,�1|�o(��sîI�q�Wr�'�d��f��D(c[e)Vx#���;��Aa������p�ns�2#��8`��m�͒�V��9�U�:R%������e�5�4����B��J-�ص��,�	h{z�U��)���N\N���֐H��Ei�\]eӆ(!Ie[��!j5�h�����*ig1�1�H ;�]a2�>	��x%1�n�HT��f(��
�RD�9�e��Ӵ�qo�w��3�b��N��{�sLCWw�,�������q���'Ӝ=#B�{�up�<	���V0$�� �"՗ՠ��ʏ���y�&��r�AY
>�厶��_^�h0ӄh}�\ԡʟ.?�m�������*�!k1����1�s·���!���,d�e�qJ��嫖?�w��mun����߈�הl �G`8�e��)vp�a��.�4���ޖi��pG�qF�)l��^��$�\3�0|Zv���l.nv+��
{�\���O�����WT��R�Q>�p��Uq�}��/����j��&�<��/,}3�7�( ��>$/�s��3%)@NQ�C�6�u��ʍ���[�7�gM�}�9�-J��.ܹ�T!��K+�Ey�o#���]k��\:WW��w�4X�D����}SfJ��є�ٶ����u`�6���^�����rJE6 �&�����L"�C�+�.��0����&cZ��dz�0%V�0` ���|&
�݊�R�Ka,���|y�oܓR�Nkc^W�D�lhg��s�9LúHH,�!f�L�Z�=�YϚ�|�BȰ>���,��M�ׯ)�xx,����K��Sź��m�<a��N�ɗm��z>���M{���	��oN n�\�}���{ysI��V�K%��9f�D��N���!��C���>*'�w�Ir��5�%�_Z���F��6ϡ��y*2�G���������P_#Eֱ����괝�Bv�t��K]v �)$��H��`gǲ��@+�Q�T��8�^t+������`���'���%P�3�1N��o��tȥC�䂵�M?A���0�,��CJt��d<����Kh���ݗ�#Fd����v�쿛*���󍫫������Ei���_ykʖ�.���}K
����Z����Lo�L�5ll��7�%@�!��L��S�������)�O+��c�$�`��n����xd䯄A��G-����6$@��ڎ@�d�K�E��K�`��cخ��&M+�U�����ڦ��D-lMXls�t)X��Q*>�������H���ִ��Z1|9z4ާ�|<�TaOVh
�,�����<�_�,�S��k����ˠ;��?F���K]x�c�<��u.HR���_�A���0�Z�f�c�E�
	�0��uo{�݃�U���DA��^ַ�����.�W"�&+�4�d�լ햃m��,��t��w,�/�?)�b�'t;��mx�n 6��3�<��o����'�)d�]�~��Cs
���m<�ϒC�� �A�r>H���)�/D�l2Y�����q��g��F��I�P�Cm.�B~B9��%9���s���Pes�3I������LOlq�Q�w�vs{/b���>�e-��4(gF���U��f⣨$B�$��e#��''Z�i��-"���Ե�%F��_�ı�XJ6@E��pz��fvH��D�U�ޑ6�K�7s\_y�`V)����F�Hr�-n�VMa�0��5덭t�y�۶��`���3��@/lbϠy�O�	Z ���kxپC��C�^��7a1�\��)�����:�����{&ᶯ��l	�B�/4 r�����,�A[�tΔ��y�- ëЩ��*H�}�EΙ�g��}�z���+���'�/s�X��t���0�>fgl�q����ݛ)�mR�.f���%���8�"����Hu �V�~��	l��T,�4K4g_���]�bU£s2��P�Dތ�N��dA�+��7�1�#yq��M�N��2�1]����������@nb��Z���w��q:;�m�>�2���7�����8�����j}<#�.�pWW�x���b�[hjD�J�n8�Y��dE-o�V,��#GtB��a�zP��K!�����Q��js
�,��$�K�ڵ:�t����x��Ws&<�4=���o���<����H���nT�h�*p�w�w���	��Jn�[Fy���f
�*S9P��*����G��J� �l�+(?Q�}��o��r���+5������[p	�Z�9�ӟ��To�.�����nvR���×iĖ��،�)�����^*v�6��.���h��/.(��g$d?��j���b&�m�"��C��Fj���#^�nm/Zg+�Lu��W��ij@�ؔc�Tv�ㅁСBU��������]�_����������V�|o�&q�{7^�"�s$�<��ڨ8�Kce��]��Sx����,�9w�m�����O�����~>�dc�n�%&���J��z�"�����y�<�'���M֖؁�S��ϻ�.����3�|�7$H+������:�+/���WUe��z����e}�!�@ͲO
:5��Ҧ����N��S��\�rD�}o���Oï��j�>��M~S����أs�k�4�c�`��lc�^�b�oά�pxpݏ��9��&�$�3~�^f����9�T*g ��Y�۶#�����_��oǍ����}0
��C�����7쀴j���k�.Þe��'q���b��ͮ�b7�_�0����)ҙT��P��y�����$�x�����!`�>�MlJ��Dv�\��H��1�ylz�iL�Su�cx�3iL;/�oO�M l}:�%}?�i h���<I�ն�d?�퀩y ��/u����R9cP���3C���8鏲��C�0<d�˓ᥭ�]�t;�F�e�'����\~	�:
2EiU�q���W���32q�����?O����UcM�8���&�X�p��i�L�J����=����lwL�_%*�tIii� �mƒ�9��lv5Kx4_�0YZLx{���h�_�tӭ�}�t|�W7bpX@$of�2�?懞��X����]͏Z�yh;��4GW@�_XE����Ҡ�ަ��OX�qÈ�����6�wAv6�������v���s4������?dcՓ�{�U�.Y�R����Ʀͣ)7A�A�"ؙ��O�I0='�Yi��>p�ɾd�+����;���4���ex�����j�aAv���}�(���uL�<��o�ZH�F�D-N�G����G���X�Xy.���5*1������쇉*yu"8{%��I�cV�a�%�D�Lb���"mz�m�#jPR���0{������Z�e�Ɓ�&�QTvL������j�kL�}���A���ӌ��S�T�����:���B��|W�FBEmX�)��dn�����dȴcT���T�	L�j�1�`FR�#m�Y���1�BϷ%�ܨ�S���<�h�迃ᦫ���ֱ!X5��g��x �KQi1&)f�v=$���J�N���Ď�W1VuJ�m!K�&��㟿��%�����E��P+��<��ڶ;�S��QQK�R�����yFQ�x  K�k[:�*�8&�a���lۋ3U�3m)9]g����XB�1YSh���ݶ'O�i�/��.���
��
�E�xn��-RpB{
D�\��J��.�b�&��I�Bpun�jIr�����􍕴0+98�&��L��/S�������bT��
�vh��+�b��-7#x��^���b�F�&�n+�J-���=���m��/��P��q������Ǹ�.�Z��~AMRse�+�JV��<q����6U\BO|��WG'X�Z!�0m�!�W4�T�T��J��86�72�n�u����*�E=�e勠��i��kmd�iy���-�����Tg��\v�v7��~T�E-�#�o:�N\��3i!R0�/�;��pI�e�N)�/Q_rvsx�K�Op����5��8�b~�:M�щqmh��$��p�A�pƹEpG�Of֔��U��%��}ϥ�}�9�H/����D���~�)�C�Sl��ǫ��?V+|E)��ُ&�n;h|u�o]?��KC�K�c<��l�[Q�x�y��|ρ}`΂0o��D,,���v�7���8����߷ ���4����,��'.Z�ވ��(� � ŷ?�@d�ǲ'�vK��?�73{?��B(�pC$fLDࡃX�0�d7p/	�3/�G"�����r�O��yi�0���MmSM�Έ������.SON���&��v��Ѭ�I�'T4��[��}L�F�aG��VB�L<նS;�hM9OP.�X��bu+��T+�$��zu�X{��6s+��'��P:�����ޜ����~yŌ'9r0굷�!�9����hB/)�RZ"���/WuZa�&6��L�4a187�m'}u�E¸-�'[���[6:�*�8�F��eq(�i�a��\�	<�l�3�  x��,��q�xe�"]��Qg3s7��s*,�G���%�+̯�$ѳ�i���*��4���Z [Pʿ۪��&�V_�F�'�F&�/��0oM�..�fy 
�������7�>J(�lj�.�r���~�J0$��mE��S��ow+BE�*�D��m.���yѮcj�V�f�x�1r����w��2A)��i���ƕ,����0T�����~ҁ�\1۝i����Z.F����I
/ɋj<=�wLVGX���P�^B�ʄ�Q��\P�U6V(,�
�_J�]*�,T��uCˊf� v�C�7�Ԑ��{W�I���ɇG]�a��W��^�'+�tSؠM�dE����S�����q4aN��.I�;"`,�k���%�c��b��mA �b�h6�kJ���<k�M+���������H�`P
 �E&��R��P��\���B* �.V�|:=$��rc��>
?nn#�>	=����Q)T�)��6/�E��=��c5���ּP1�=���)�!%��H�&�@�ַ�N��dZ��)&�j��Uᆂ�!�'�"{%F#L(�n&S�s_�A"@�����4A���6��䳣��9}�ϱׅ��z�}FJۧ��������&I$
�oz[�����S���)���/�4���U\_�!=vu��KKpr+L1)):� ��z�iz�2C�q��|v(�)Cv[p5�4/iaۋ��g�'��~�>��O�ǽ&�������]
�T�Ր�	Y��ZDM��uǜ.�M��������Q�_g�ň����ͭ�ػ2Ւ�o�A��kX:�#%w�e�C�=�7ͫN�̏�h#~��
�
?BZ
9�+m3{���l���7���/EX�q��i�ʿ��t�(�Vu]�~4q|�ӓ��H%H&4f���������R�)JF��g�C�? �97���$��Ա��Q���?���Ui
� ���+^;� T�tp�)]����Xu�9��n�l��=�ΰ.�w�����qS��@o�¹i��1��H`������lT0k�!Iv�i��C���r�sPo�we.l�䇶�3�a��4mS7Ұ
�[�i�3Oj��~��U����n\@|�qQ�����(8��=_�8��(���.�/I�⃑LE���{��R��s�lI �������"%����ͭ.&�s,$�|����q��-]�<%B|����b3͡��$Ԏ�#�oQ'�e�K�Ƀ���j&�z���&�2�zSzGf��	�"�1KE}���2Ѝ07�+,T��̷�%%y�L����V��?�v�b��e��T�O�R��q��%��[����E9_j�?4��ww��>S�}�uۖ��~��`/�����.Vj�{64g�ū55�M����� 0i�<��
�S�vn����R ���R�K���R��d�C�:�d��� >*K�ձ,4ʩ��C�ek).QZ1�(�2��*��t����u��e�(��U} ��}d��:B(O���D����J8Q٧�zL�C�|p/�'[D�ׂ���y9Z���/���n��l-Z�&o.��W�� �EA�D!�ĤJ�l)�8�Y���˴9�,8L�ʼ�1�q1��ѝ�����) W���92��'�U�Wx�q��Q����P.�9 ?z��WO U�N��73#8}��@��z`����A�)����C�n����g���� ^�k:��@J�	s��-�gQ�zz��mF�K���DYa?��A���R��v��A��K�!�!�9=��&`<��>��M�8�~7U6��H�玕���M���~O�Ѝ��-��ۛ������J�=�H(��B�*���}`�_A�M����b��ޣVۭ}��U�=e��0�5�A�OB�#�ʖbY�r6�m/�������ZI��;]u�Xd��$V=�-��o�Ӂ�R�H ���A�) �����M�0�-7 �I�t����2�k7H��䎊�#�pr_$���ڄc��,	|��NA��k�G��)�k>[�������88gdiR��9��ވ�U�a.R��딛�ꁶP��٢~׀�����ծ+=��ÏjF>:IװE�a?��y��]`�����e��*�d�,�\7�®�j̖�ɡ���K�#q���i�M\r����#n���錄1�뚉��TM�"�f��t���}׮\��r�A>CD��=�ǚ�\�]����d��->�lq$j3��c�Y#�A-������%H�,��H��*��? ���4g���pTӷ��r:�_�Uz��b��e0�H˛m��I�~֚�f�rĂ�ݒI#�k7bH11
P*�.3�|*ѥiy$Vz��ga��Jg���݇��@�Ƴ{�PH{�ܶ�m\���׏ h�1	[�eH�#�Jq� B#�`P|�-�1��f�����ToW��hMY?-��~���էd�K��6ѐUL��.R�5�'�"IQg5g�~��G�"f)ݶ:���N2Z�|����_����F7ZN�	�=�u�f��?}�P��ѼO8�f�Η�8c� Cf~�Y;�D����{�G��@�b� j�H���q��/^��zl]�uP��s����\��<��m&�'���*��L�,�i�]�M~��+D)��Q������Eѻޱ;X_r|�����5��CҼf{pSe~ǧ�CO�h+M���M"�5J����]���w���p��c��Z�̚��D��8V1[W-|���~N�.���t��Wا.旈���@�t�����G�0�<ba���=�d~�d	r�`Q�R�ff��,�kr��FEH�hvjV�>�u^��w;*���h���W�z	ϫ��~v1�����Y�m7�U���88���q-�Ou#G�[[;��Ĉ���2�\,g�O��g�������(�U��4?ٍ����d���{��FF��r6���@ l��(��we�����]ط�/����F��Ҏ�$E'�9�!"5	NP���=3V˳&"曇�]�x窚��O�Ù��H��2�e48s2���3�����.�Ma�%FT�0�zjg;+Q�����OHHKa̾��x�8<��=��3��_9-��nx�@F����`X;`" �Z�
�OO��؏@��I/P��>J������i����zЅ�
-��=��sr,�s2�m�r��V܎R��W�x�9	i�^�Ε>d
EI�sh 1�y��FҨ���L�\���e)b�0EY�Y�~*t�d�@sh{�"��z�H����L
[�R��� G	ͦ���=*{T|��~0*�+ ��*QO�>��5�J�����b�gA+8�Ε�n�(8�#�g[�o�H
�.�!�ų� aD資'�}�a�9
j�$��6[Il'�xN��|+p}�:J�B�[⇚]��p>���'!A=d�8ܒ���3-� �R�Y�������A�!O�gg�G�A|=AV0�rx���wl��
���I�X��r��>*�y�dٌˇ!�6��9��!K&��Bv��ci6�u�}��9� �T�w��;�1&5ǵs?>���]Pt��t&'r���Hf:K���Mfu
E��WC��$�&R �D-ڢN�5ڃ����ٗ���=���%��H�a+?������f�?��}P@S��s3`X�'�����*߀VH�����Ԋ�I8���o�����ڰ�U�
�u�����~��6�#p�{���ɀ��!�t�/2�);�o���8�;�A	��LQ乓�,�>����	o���)���r���f2��c��h � er$��D�Vp��|4W�e 3k�F�����������U)��֘�����ۆ�DE����'�J6�"��@�)�֩�2#�@4ʢ錭xvgKr��<?�7O0o�^<����R�F4</�a�w��� ��?��f��L̅���"�[T�@���z[�<�3jQ�����&�qu�	��*�u���?���u,��x��]���R��}��xE�o�iˋ���ԯ���
J���X8�Ԯ-KyB�	�����a@I�s���^�����-ɥY,v�|�:cg�%��*�tǕLkycE�~*�����?����c*I'�w����g& ��:,�t^��+gf����6����'T	Hru�p!��&�lӰ��0*�3{m����k�^�}� �����n8sJ2C���ot~����=��"�NUtI�GC;�DCs�8f�t<�$ e���t�rWu������ѣ���6����Я4���Bq�U��8�t\�O뮡+@U��v/�7�\�7��Q.��0NA�W�ǆ���I�x�D���t�T�ч1�����ұ�2�/����=iͱ��������?f4���;���g�� �J�F�6H����zXX0i���5gN��~ڀ�D��0O��K�o�,��Y��}�s��SU�#�ش'pJ��Vf⇨��@"����>���m�N���g�K���k�����˥��WQ9#������c"߸}�7��^]d��N\���'�< ���|����q�#u�4k� �#J;&y�K�Z�-~���t�%[�%�(�T+��ʓk,A�p^�@&��0�0�/�M�+jQ�usbwB�ͭq�7���p���ju�m}�z��Aq�_By&d��nr��ɳ�F,��A�Y�N�{�L,:�6�o�Ig˷8���a��j��7�������s�>s�S$>�u|rGȩC��m��3^�L�Ò�Y�YY~�ޤj>3p���"ϛ��(b�BRPk+p�\��4X�ڬ�m��t�v@Ox�ւO���ٽ�"�Ս/��k�!����|��.�bV��0Z:9ZpZ?�a3k���G��ߞ�q0=�չ��R�g6_N6ae������owR(mt���$ϼ(E�ك���,��g��[P8�����֝�a,���j��'�x�R�4�`�5k\��g>������R��7N��l]�W�$_^���.̎O��j<�!c(>zb��/�|�Y��Զy�/��*���T�_�o�(�|F����K|�7���=��/�����*����٧�.P��)��������͔N>V�O����K.�WS����Tx���������K�:��p3e�k�
8���а�k'��)�Y�	ͱ%urdq�qU)y�^f�9���wXn*e!�4d�<�2�wy|�Z��nEAjX�;�0��~"�ì�i,�w�,X�HIw�2�#?�&U��dE�f�)uy��#jz�Q
�8�-M�@����~�4�1-m��:�������~�o� O���8
��5�FT�%�!�~��$v��\�k^��!'�����y�ȣ��1c~!��
VRY�ǉ���
�?��NeA�dg�:u�К���2.�`�U�kj$�i� ��D!orʂ�b��Xw�\o>�!AV�4$F�d�%��F����L�H�
���;��a�^�u7��L�N�Q7��_	�l��/�ǅ�\ˁ��5qIl˒��Y?�{�G�1d�	,�f��g�d�[K�ڰp�դY+w�F«��U_�hu��'��9����S82���"\VøpJ��m�~{l�x1O��$����F��TXRS�y`4��qH�f<N�Ԝ8��F3һd3�������\R�*�%�H6M��u����蠻o[����y��o���(��r�rGl(�\2� ƌ�*�z���M%��Jo6�@hWD��+���k�ㆶ+WNtJ��\QX����3�<X�{���4R�O���MzM�P�K)H���6�2��̈���{��`�S�3��&�_�=��'ʧ�g�Z2�+���:���T|kv�4�#X8HMi��4ϭ�5D.�L� S#ߙ�՜Pg(&�����x��E23f��N4���;\��,��+��s��`�8UH���u��0Y�+���;���C�|��i&/����Rdw�=�X}�>���~���& ���B���
X�����F�9UxJ�9"�+���@��{��X�@�+��>�K^��*b7TU��MH��4�6����{r[ub/Zcd���"گ���i=��g1����\ל�y�02�j4��j��+ʄ� @h�ҵʺ�Qu�G�*����\+bOo5���٢���>��jY����!�Q'�t��O�Xw����!�5@f5�	�R�!��� b7���M�������ҕb�1X��_��w����-{�[<��˅#u�]=#��[T���i>9�p��3j���Q�qm��Gؒ��Ӕ2A&	�E7�d��@?Sqo\��[�An9�τ�D0�?��Oh;�鸓��/4c�5���W��^�iW��U����#ud�eXq\c�Ɛ��W��qI8�4߻G����P��a�����x~��[�q�b/J�7���;�_wT{E~��;ЛX�]�[�P?�֌��m,�|�Nk��3�I����=���Ҡ�5T��03x쓫����$[��Ѱ�)��^�,���Y�C�b;��)��'oҋ!Kr���lX�"x�s��Ϛ:f|'|<g��v`�%,<"��ܛpm�O6��V
)��.���҄�Zk�ȹ� �*�D��3�T�B�g���ߤ>X�[+�pS}��u��O
�☴ԴM�����^��e�{O�.�:���w�Ee�:�yN�=���.O��d�dFޟ��t��F`������c5�m��/`S�j!m���,�
��k�O�D=d@�pp��ޖ�1L��.;�k��x��R��G3��3�S����z6��o��WU�c
���F?ix�B<f$��*F.��-=@8j�q����n\;d�Y��Ü��=ثߠ����#���{��	/��Z�S���t�x��ǘ�� �7,[]�g-G���tȷ����P��1ٯ�*Ō)���|�R�a�&O��ܳ|kc�)G���q=(��hfCD{!2��@{��w
�Ə�lblz�O)��Ң�c����,RQ��Ξ$-D1c��PފT�+�e�:�^ɑ>U�~;Ն=+�W��`\��JeҸ��6�)�MSp#����Fl���~��kavY,N��pg�98*�5��*서�x�ږ1��D/h�xn��������9j�^GT⹞���%���zQ6k�4����#�E�����`��}y<<ќú�C��0�f��B�oD��)J3̈y^~�EΘ,��j��!{�T,yhltԗ�pBG�U�논�y���=���Pı�z�^��H��o�+����5�����{p8l�ߚ�R�I��Bh�J^��0�6\����9E�{�(�Άpې��;����G|a�E��������;�(wO�լK&+Y���:ؗ'3�~3I��z2ƣ|�v6�+O=�$@�,).�;�&��O�F�*Rz�7I��P:>��c->�P��^TF��6�!��
1�U��Y_�J�=���F3���`�9J��']�S�Ѧ��.l�"����� �ny���<���F����%b�U>�<T�.��D3PE�^P8M���2�!h�`J�փ�*;��
���0b]��_U����Z����d�Iz�zSHȆ�\��6��H��6�sfqO'���3���J֮�������y'9:A�ؔ���X���_�r�^��B�#���V����p9j�����+GǇ��D�He�����{�eiU"�y���']u�]ܓ��\���b���@I0����Dq�ñ�U*눖73��x$�rp��)Χ��"����H�n�����
��hɰP!���ƕF
���L�`<G,ꛆ3����i�E_�〘D�Ɛ4!��ϝ��Nf�9+��F��%�>�1�b$N��*���$\�pA������: 8*.7S�$ea�S	���V���]S*� V�T2ɻ�c:�h�!3g"&��RQ��5�"Y���)/Y�}�_��?��ݨ��|�Wr����0㼦�����ٶv�'�1s�yEf_�+�p.� ��M�P����9�}lu�Bۼ\a�.��B0�� ܁ o#�vF���f,@j��D��3c�>�\	�l`R9��G�S���?��f����:Z���l�hw�Zk]�e���C���:�tRg���i�!��K��q��1�)����A�Ih�{+�L�zB�.`ޙ�p& Q�
C�b�k2�'b���
��46��q����v�wˀiпR�k�?�K3n�9�{߄��5, ��W�ooɥ>���z|�'p��>7D5L�]�4ҥorA�:	A��'�wCi�o����_XdR�
hh{wCJ�U��7*�I|-P��YY�~�T]1�ե���4�>.W�<�Z���Z�iQ�aB�ʴ�t�!�q����'�j���΅%�����F���0�)�+��d1����=��{󾺩��|���9����!%t`���9��,q K�ؒr�9���	�%
��'$yF Xc����#P�JR���)7�B�K�<���<Π���IBq�2�?����������4��1�r��#����8Yh[ު�j�6���S(��*�W�'sI��Q`�����TN!��p��	�H+�*���h��$7���'*�<%�#��ax�gQ�Zݟ^G?#�a����A�zo�n�*���(��k�:*AzŪMÄ*&�Î+������L�7�PY����ދŬ�S��)션�;���(��:��#�{�����<�2�;BE��|���Fĩ��}���U�<FoW���k{��{z��!$g��l��G��.o�Ҵ���\_��N����\�I}Av���I��gh�#Òn�0pW]\u[]zUב��ո�L��Sc�o��n����8��Y^Bt^�X69�PY���Ԫ���Q��K�[�I�+/N���>�X��~�m�x
V�����달Q�1�X%O�ddZC�J�1p6E�M�����^dX-��hI�'���Xx�,�4�9�&_���4ײ���D�j��W�u ����U]���X�v�:kj�=D���Rei�i�������o'�̫R'斧��P���✁Y�x��E ��
R�Ԕ7g���=Ձe;��ȭ�i������b�`Y�d��Ec�?\i�6�CDc���k�1'9�Z ȉ��(��b!D�Q � h�T.֏���̝qǒ<
�����.~_��
 p��/1��W��>� �1��S��� XtZ���R�}7N�~��Z�H)��b2�˷h�$�@�� 	_;���҈�޼<�t���l�b>P��Yzp�����g���2H���D��_�'��|YwcY7e��r�Oec�"ޤ���-S1NǱ��w�yݡ��*��kG����ƅ�ؤ�<8:�i�7Y���֦���Z]LjΜ���DO3��w۞]�����nY��wHvl��~�c�w��K`�JZ]ʃ@�]N5��8��4%�7��J�&\]�<�
��g�8R�"�A�~V��$Z���q�a�6�(��H�@���9��ZA�R���Ć_�N�����`��6��v���f���L��̱ē�x�C>�`�P{����{�Q�=1��D��K�z�PY7^.�^��!�?��i�dA衲���+������s$��Q��ˈёh�l�i_�,F�#}`������Hh�:@Q�ӝ���}Z���/B^��?�e�ͯ#��ٌ1��fߩecZ^�AR|��q1)�b5�H���?���)��7�Z L�G�(l8��ٓĩ��is��Ij� �+`��������eSn��52�[F��q2U�!2����S����Vg�m�-<���%���O�s�Yf�T&��2�c�[��k���u�S��n0x>[I�*﷮�U�pW5��߈�N0�;��"�0�~�F�H���G��cI��4i�Τ�r�~�QI9)�'9SU#�s^ą#��Q�P|�z�C�άC��k����/_z%mH��s]�C�-]�����Q^�bda+^��Q�+�7�d*�oZ�B:���ކ<^S�J�ݷ���������/��3/���q�X\��3�v�C/'��v��T�F���>�Vou�*������/�:`���t�/�dw� x�ɘE㞣��E���A��b�Q���+m�E}�]5���cc�%c�Z�M��� �a������,����ʌȪz��_�l xI�h3�?���!�uVk��}�?6Kks��yOb�	-�����@��V����%���&�� })�������|�Q��\U(�h%ם�9O�J�]�#�b�(�t��xg�#�+CP%/��v�6�
��oo���A�bdD�Q?�T&@3Y��Eغ,_�R��KЙ��b �W(��mL�1f�I�b���J�3�ά�J�5>����?���OQ!^�� ��	Dg���9"
���jn@��C�w^oaԊ�'��R�߽]W��,��;r��`�@�vRBdI�Eqn��>G�
�"ش&��E"���(�^���L�L���}����f�U�u���ވrzY���e�{��vK�O��j����D��TV�7劷hQa�|] �X+؉I?`c�X��v��g�x�0©��=��3�ۥu�}����~w׃A����&��*��5F�@�OL��,� ����gءʇ�F�lq,��ivr���{�r�����H��ᙰ-'<y�p�}r��rI+z-z��`SX,\\���]����q��+R�4�`��{]|׺=��\d<j�z&�E�����v�7h�4��+v.Ԙ��#m�!�4��T3M���KN��<��Pk��;���g�EwR�j�������N�ty��՟�t�L�5�'�!��4*q�'~�۳�|�V�ؘ�	����C�w�{��6{iC�%b���xd��A��Ra����(��q�Je��PvQy�j3�x���P��!A*u��Ǒa�����<l%,c�Ŵ ���,����2Њ$)w2���l.Fcn�&�����8��;�����|؂oBXs
�A=��?�9���I�ӛ���@����F_��;�!ҘX��j|�F��,!�X(��ڝB���;��l�_�x��q��@�kF���HXf�� ���"I�(ڹ,�ܞ1�n����}$�0"�2�7J<�-�	{r&�^�����w�<��-��L0��Ռ�c�-��[4R������Yky-K�p�Z�	�Y�S��/=Gr��}���͆m�m:�X�ᮩ_\��P]*{��U��;L%�s��x����<N3���w��Z�a��RS�hI�WI�L���X���Z`B��.�?��uo�s�&���~��vPڷ�F*�*��Q{߉vrV��rK��V~Or_�p��=,��#hε,��}��}�<?�ɗC��b�Z�8�]N��KI��m�u����>����Z��C��<�:籧m�3�?����` 9�鷝�5���.�%Pu�i��z��}�J(�N3���+�Ёpv��3�����	ߛ�@)����,�g��cG�'z �����Gft���	v�Ԡ���}A~d�n"N��7!WnL�P{�����{�<�df����1;��!;a@��/��y��O^uR*�KX��Ӟ��%��ք&��_��A���fVf��m���??�79+�j�Y�Ui�)#ώ��)z��ϋ$$B÷B4=�b���9�;���:�i������D������3Jx�R����T��_Pc-Uot6�t�h����?*�~e�ն@(��D�j/ X�g��t�������"�wވɧ��S���SEP����@��|� ���E���t�ةt�`׳����h�s5�j��ߢ��zG�iӒ~��I�q��бKc,^�c��;�jf��Mpx|��"%۽�2u5. $�p���:�5Ew␊��;������1��ٰ$�:퇔����e�h�UQ�J���<J|��'n�[�rr�7�Fcυ��&c�\~�n}�!�\���7�����dK��T�HW;�������U?��{⚌&/����=Q�UN��z���nN���Oh`�+���,��℗�j>�������)o7@���]��Ǖ�,t� ��>2;0&\n(89�!��$%&iT
�nB'X�pFѻ �x��Њ�Ԉ�Ӛ	u�
���t�uؔ�� 8�����ěd�X�k`�v����uJTAbA	b
u��B.ME��SwE�8}lS	�ީ����5h��`0ZNp�/g� �:`�4��B
ަ�`8�{����`�Qǭ�D��9q�?�p8N�&�d@�jn��W����񱲽��^�(y[�������*>���gg�J�������Ȫ΍���:�;��Ed�?u�����H`P��A�Iڰt��"��xyU
[��_�N��(��(㶽�@^����<쫁�5AD͎~�[ʃl��ß��]�g�pH/��ٞO�:��{ͨ���`NCʍ�uyW�,��U<��n�wP�j�xrER�W`�x��̈́*�T�BY�
��9�˅�`jB�֠9�ׅii�ؿVm�}���h�[�p���x� g�f����Y�c�>8�nĀ<�E���w0d�e_a��X��b�r.�EP� �}�pqx���v����D��М�@�h�lWK�颈�R�m�oYzw"V�)�+d5��fG}y
3X�'�݉,�W��	QD�7u�&EB֗�e��,I��YMpj��t:�a]~vPyLN��Zݐ�P�z8���p���Y�b՞,�?��,ս� X��
2��!�Յ��_��m���~Y�y�����	N.�J7��?���M�Mk�\+s[���1�ȿ8��b�i$�R؟&d�h]�{�:v\v*�q�����GSϤ�jW��B�R'�Y2`�v�V����_�/?�Ձ}P,�7\�c>�E��w�;�~���?�w��~짣Z'V�gS�Ѝ`+���d�~�%�)Ǉ	�r��=�˱ot��cyE6i�uȿ������oY�f,�Q�/ˇ,)��̄�0c����XG��	ܹQ�<B&r��ڢ��n��N%Y������!MLPW#	3���k6�'9;�+2�;�?m��냏D��V>��U�N���ykm<�����������sFnJ���2]]���z��!��cj�� ������7����^ Mg@��T5�wt%�Az��Z���)�Yd%s�}4�r��mq6C~-Ұ&w�[���!�p���s��a!?%9>`���~רD�W
�[�0�W>t,�sR�i(c���[��#IT+�[�z
p��u��XTr�.׭ظ��N1&��>��3	?�;y���S0�/Oɗ!B����.t�y�<' I��ɠ�q��%�3|�jaJ�LQ�i��I�c3<��C���  <��rP1��*�HT�MH�[Ɲ���Щ����f\�*7ɭ[�лQ��N����q][�,�׼������H�'8�i���+�����	��$Lޣ�3a0/X���輗�t6$���Z������̹h��:��Ɠɾ{?�^{�e~g�Y����wD���2i�nψ� ����\4������:���A�r�BG+�(�Y�h�&EhY���G|�F���Vq�5���.���=s򙝈��&�>"1��A�p gˇ��U{��<A�@�B�c�sX��O��~1�w65����	%ZM߈���_��%c_Z��̷rWz0�L׉�hʹ����������F�{g-�3��������NACUEn�t��B^"m��,����A8�t���^w4��u���;훀d��C�k%��ԯ�/�6�cƎ���lV�EJ���0=��/1`&�K1���$�y��-Rb�m�����eD1" �Xo��o���q���eR��_|�	[?2�P�D�o$3b4�D�g�k�!K�5�*����0�|EQN\$V��5p�T�Qg�����M�U����5���Dy���j�#ݵ�f�kF䬣~ ����t+�/�Gc�+;�^�s�͉*��)��,�'Q�o�,��E�g�ү"_�=q���{�O$Uԇ"����Q����n�Ξw۫4@=���$��]� �mG���C��b��E/i�?�'?UT:)M�%���\՜>H���Ǯ�~�P>�n�шz�'Q���p���"�N�1��/�����+�a�p�����8Y8VhE49�������ag��u���aKDs���������˝t�M��Ao�����R���"��<���:�����D9�g�1�S�2�Lw����,z�? W��v����puDǄ������,c�7�t���"��!܌ԯ�-��bu�V"q9l#q���3��ў��K���J�nC���-)q�~����$#%�c��Wq
Y�ൔ)9жr96-���6G�1)2� {t�N���a<�Nvq�0f�SB�L�Rs�s�.��>��~L����9�clt�Ug���(����#ئ8�3N~ݸ����PL(8w�\f	�CZ�_>���,��ە�6d6b��L v��0a�-A[B�#5�_���G⻟I.��B�`a6?>����Pl�!C���2]�����00����,����RJ�Q�Cm��a��/���\�zP:��N���{�ꞽ���\�����Z)F�\���+�8�2�Oؾ���+M�#�R%�9���0/�\�Vy�Z��*��l&��RTMj�SU���q?�fը��7]��2B�� ~o����ަ�b�����āͭӃ?ڂY�]��J8?�E��vI-� 	6��/9���#��Ohp��+6�I9dp����*_sWR��W>�PCp�݃�Z�� �m�@��M����mv/P���2�!̭��`�cxUQ�Ͱ���1;�]L����^���l�	[�pa ����c�	z�ۋ�뀥B�X�K�`#�d�b�V��m�b����-tgY��d��b,�IC'�G�D$4��1 #�ͫ�l�1d���|���yz�4�7�?'UqnV�
��V�Uf4@��U��a�=���W�8���蟝�U����X�1��g-.H,���ߛ�<�J,����8�F�u�{�����sJ�ˮ��6 L�č7u��'�==��Jag�g�2Jt#px�L��)?P<y/ ӽ�����5���=n�0�����<o�n��`��eV�{=%���z��;q�Y䩴���U��k�KZ�t��FBd:�B�R��z�o�G#���%��Cn���S� ��ߑt���M��%�ѣ�Ϙ��kh���Pn3��W��d�}At��? "	]C�1"��ʮx7�E�F�Gpy���t���q�US��0�-"������dc���,��On����M��J�1�3��CI�����I[~*%ϒ�s��僆s![k�Ų8�:q�5�qt25f���U�в6��� 	�5�6}���~�����;�x����.��2�޻�d�Gĝ{{Е��,����47�ے���l��8�BK���c�����LڹW�0���[�۬1oʮ+$��cΈ�O)�7��W��>R��Ԋ�jUYq�V, !��p��3*�Lb��O��ݟ���=D��6fm����(��|����1l�Ta,��R�M����&�g�!g�>|������ijS��AK��g�.B8���~��`�@_��PB�N^�OzL��\��@䚾��)�R�N���ʨ��+r��CLO�P��/���ڑ���Sr�y�4�����Z[��I���7�Ҋ�.TcW��
T�@�"J8Y7KhX�fi(u��*�`qW*8�!`F1�-R��ў0Ϝ@b8E��`���q8���%��v��vb�@��y�b��/;qPց^}��媢!�3���	�0��8����"���G�Q[qhl3�J�_�%�Y%���M
*����Zw�S�����.`�F50�+��%5{��rY�<[QK���U��W8]󘺎��H,��<o���-�9ة�	�㡳�E�3��|�i�<����&^S����wl���7o��P̼�8��������S�ɽ��[E�!_��2�q�����?J4�<�;79��o�'./��S��Jo�w5�����\�,����]`����.��ڻ43�Yb�m�%�0 3Kj��d�;���a�"�i��i�x�q�}�������<O5&�=�6��z�ujk����/����W����v�Z_~��]�@�GYU1 z@�X��PÇu���0_�/lA�L,�E�C���Q��f.+�2[�-`v������?���A~=�{����]��H�bxnVq�P���1����ܕ�?g��B?�U���w��~-,l-Lb�X`�`�f��DEĠ��	���eU�Hꭜ�o�:F ��ƃd�"�#/�q����������`ɩ���'H�����Ma�q����L��E�+��%9RF��O25Lk/�TO5s�ExJ))�P;��	7M3�~�I��S99Ϭm.m�}9b�� ��0��H��z=���(!�;�T�4 LT<��[��1."��c�[G�=��7��QT�J�i���M]�G�?� ����[ %�e�YYvM�Ug�ľ��ps1�ˆ�(����]٭!�:��&\o!��S(��Ro�6Ex��O筺R����V{'|�ܽ-aBŝ�]r�������"5�p����n� ����9�cu����n@P��=�i��_3��z�mf5(�S��a_�'%���%TO���=��Z��&�F( ���#D^���{�K�2������!s���ѱ�w!.f�S�G�\%p����Zf)�=i������0��׺�j�e"'�#ghH?L��g"'�&�.���^��9A�W��J�ў3����R�I�N�n!o,��ɽ��D����cy#���j�sC����6����*i�G�5�2�+�6�UB����8��"^L��3j�31�or�5��E��Z����w�����~[�~��_��=	���<��%�C>��7�u���Q}b��oA�pS��e�%@�����8]�d�垩L ����(i-{d3�D��ї��D>��M������$����S?�+Y�~�d�K��Oq/�vcE���;��q,卧"��U�gz}���⡤��Ye�Ã�#f�__�d6u�	�˻w�1\���Y.Q�Ro�UL�A��hy�&�-�%��ꖠvK���o��=jk)>�'���d�P���U�+���d*��a}t��	�'0��X���<7"í���Z�č�������ڬ��;�s�|`���z��?��e
�`��l�+�!��'�������/�"��h����$��A��2�f��]}��ȓ'/��TI\W�059�N������Xr	��E�����P�]د�r5�5&$i�d6	�3�5a�@���Ȅݰ#��ձ^�iX_�;)o9%~���<�}lZyqj�-�u�L^���7�C��^:)r��b�#��� 1��O�z��d*�DRq��ܤ����?��ΰ�^�qf~yrC�?p��Lh�hȇģ�܉�����)<�sw��8B%���-zd�f9�NInR<Z��G���}�Ȱ�_�^��Fd�|��3���c?= f� ~!TJ��J�i��4Z�W->�4���3ԝy���-?l��OH�K�o�*=�jJ��tK�ؠ��F��Z�R�%����׹�ea���:�eV�l9�a�J�e����!�/��,V��y/wHn�7ھ:����ߪ5�e���'tٚE?��n9\�4CXBD���bM���b"8 ���C.���үk�y�7î9>w�*�w�������rE��)f(C,B�ǆ6�*��7	'�]�&�"�����n�����_H���t@�-���q����傩��V�+d~s�Do�(�2��}q���i�#�֭t;��b��KJu���S�kOP��u���|��y�Q։L�ܸ���r����М$�&��ۇ�C8_G:��3s��(��&sjE��ʦ�R ���~�i���yŇ�������zv���B�.T�����y�H&�ʹ�Zv%F=W����2. �n���:�+uw�\M��C7���ݨ��AS��;Kk ^@[�f����I��A�%=xe��r��o8�n7" İVN�c��y��*z���GM��ה&��S�2�����d��0�j�Σ���A/���i�`?w�~���O�<�+����f$^8��ZűY��1n*�B��L����m�<��	H�T�jo	�y\�Ǝw�a~�K�rB�!�D�8��}���+O���]����TnBdt�{�����\MupiP�"��:�@!A��l�8��ܢTǤ,���,�\�ދ=}=�%u�ݣ�$�/��׀��SK
pʰfɇ4$�1x�V��Q����#		y��z�CA��>z���dM�.-o��O�EOw����Mg%�=�
�B"A�,(d�6~��곏@��'\-�>߈a��������h|<Jy���.K2E D1��dS���nC2��.���n�^�I�S�g�#C��LY�+h��I����\5�GW�����Z��$���2n�Ώᄲ<��5����-Ӌ��W��˻�i0�x�Ya0��UL�q�S�кd>$�"���S`u��-���~��bzp�RJ�:1���Y:f��Q�	���l�Su�'A&����꬐��|B��"��6�^�?d̡���
|$�O�z7�k\���h��.�Ͷ�Ƃ����F�������NM��~6e�m�=یɣ�ڝ�e8X�o�/����ǔ'3��Q(�H��!���tiyctˤ�W(��%���'��	S��۶�E��re`7��z3ӛ�U5؃}Ϋ:B�?O�%���Fm��g��$�����'Yh�����D�e$�m�MD�{�Uϓ�����^U�]��r��JZ��hg��>B)�A�a�K��ߨ���3�e^^`����qN	|��֕~���$���� �7�b�9�Hq<��6����"i�}�nx�4��v p�_�~#�+���2������#�:�u�������)��k�� ��U�����z���@^����ݫ爋A�#O,��4�'CV?��PO��GgۉNT�3�w��a�*vtcP'!/Z!���⣱���ɇ�-���C�KHFO΄�wy?�K&!8[8�N��s��rކ��"�"�8�� E�a���`Ry�f���eW�wX��t^�k�ǎݭ֥�[�[����NL�<;�v5����4�A��)�A��um�O�t���܏p!| Yܐ���ɣO��1)�B�\�g3*en��c���˓#H��Q���'����f�k2�p��ðJYl��-���5�U�����,����^p:�uƂZX:�΋h9Ϭ�O�X�%�P��h@z�&�Ϻ������Ռ�{�VGI�&��Z	�����֏�ߎg6x��F:��+\]�j<�4"���{l!� '`R հmW��ByW��f� h�ɨ�*�����˛�݇w����HLe���]�� �l��a+{Dj�jAN\7���q66�c��ft��%>3�:ܑ��Vn4�Ĥ��᪂�")�Z�H[�� ���W���.Ł��V�Vv�� �]�IN}^�"�_1-��-_�zX`FF�&��u��@4�Hi����E�l�.�����E�߷?�i�DE�e` �+���t����<�w��o��)ؓ.�~ߩ��1;�1tI�P��W�<s7�s�:�@��ϗ9��pd4�{S���x�����ؕ�;;��a�����`kuv4��c��"��Aλ �MZ�_2���*sB�bi]������H�\�69ω͐�X|P��u�Vo5E?rr�pV'�����l?�<c[4�;;�'�nS��Gk��R�x��������Ȯ�}���%�ּ���h^p��;�arz����y���D�l�Lu�4�P�@�$kZ��D�ݒoM�M"�=B�L�4�˯�g����ɝD�?�W��$�q���MZ��	i�;�0�O�2�	f��V]�b�Ƈ4����F�Â�E-N$oR�(�E� �k{���Bx��c᠓�ܪ8��T�m�9���شY��+�pQ� ��x�-xB��;M�\r�Ύ��vܧ�6��"��]PG������k\��3J^�Y*	9�բ���1Zr�:����/���g��]�&1�c*5��(����^}�gm� �)\��9H���\ߤ Â2Q>�����SޭC�=宍���s�ɮʫ¯vk�����d3k�*�IS��`��]{��"�#�2K�d�v�ܸ_U
�Ƭ��xk�S�8���j��<{L����ŌӠ�>�y�h�6C���Dv�]�³c�=1!ږU�h�,��:is(�b���ph;'i�[4��"�_�]�S_�7���{�E���m2���
�6[K�2��)"a[H��|j�j&����'0��~�����罔��LI+�-�ɳfS����J��N����F��p��![wS0���Ѫ2�� ����3;"yT��tJT�IV��,�U��q�	}@@m�D�|�%G�$�9�>��M�'�	0S� X0���-;���Ǌ0k�ff����T����Ga�9���^�>�N��:��oAp��}CX@��98*Yhk;A�l���*�)&�q�E֗�V�*3�-`v��{$�=Y/�ٹBt�G�e�j�AT�G �/x QQ��6�q���W�����э���Mi��޹�Q;p�hֵ��.�XJƌh��ʆ��fPWi#��ȡ�� 6��2T&���\8��>����E�@�(3�h\�R�.>�r��a?�s��z��yg�����Ls�g��-�c��v���k1N�J9�?�i�x�&�7�� YV��ّY3��a'h��س{�I��p��ۂJ�7G��r�P1��f�C�K�����a:��� �6u��S��\	�;u�����J�H��*��!)��6���4=n�\�k&&��z�n��yJ�/�>�e�أ�P�b���/�t4)��F�R	꼽`M�������ѪAY�/ѩ�h��2�T�6<7��qE����J�d�\�.]���ڶ��*����r�s�u6�(3�|e�s%�h�X;�|���Hઉ�f���uQ�v�UӲHbf�1���G�F2h�I O�s��~�lmCJJH��M�`�n��,trNj�_রI���+���%
5�QhÒ&���ޭ���#��~�J�Ġ���$m��W�j����G9ꄹ�S���Xx���
��'�� �R�!�j`C������։���! 6	���H^�CuL�-�;�����?Vڎ���R.���M8t�����ʒ�D(;(?��p�R~9�Vޤ���q��޽C��$6�����In��i/�lG�l��⿒��Z�6�3�p��'�75��cV����_3�+��٩&�w��'�5��2�7�/oח�^?��� �������>��XϞ3Րfȩgs��oY�/�Cu�؍6g�V�i�W= �A�9��Ev-��>�
HZ��_��� j�B�@�婍4|����~4���|�P�7]�x�ZC�h_�^�Y�'ʔ����c��q�X�zЇ�ϛ� ���C
�ٔ����欧%�Y{��k�;�Q	�=� e���Ob�"�#*Go��MW۠���o�G,���5,����u�������MБӛȮi0Sk�����[��i��qJ/�X��!s
1\A�@o����to�5S������b� �t"�0g��:�߫ҋ�;dP�{Q��-,��)�?�+��:\i˥I��G���/����^K��
��ԭ�!�.a���_�����5�Ɏ=c򶞰s�Xs���w�H��f����v��?����>^r�Dmp����l۞���дo�wKEz8M�5/-m�K�)ޡ��O��3���U:��B���_&�%;�s�.7�����&�_�;�So&f���HM1Hɬ|������UT�	,^�I{̍�Ɔ�їH�T'(.�!�&�f��q�.�%O'&�	f��xcGW�6�h����K@D{-+��ﭝ&0&�O��(�]y>��LE� �O��7eع%�ly��`%�V o�hv��ʚl�ȕXeO�G�A���T��I�I�072P�� @�w���)	LȀס����3�d�\�2�
���{�ʈc�t/M�Ry>ϛN�7.���e�@�น_ i}��({J�8E�}{��H����~d�����z�t�h|�~# �Z�,�B4��	,N.�$�7�3�'�_��4J�h�]5�l�sFDnM�����1r�^�2�a�0�]y�寸�ּn��<�yH �B��6^6�a �� [Σy�%�����qe�xQ��g��y����r����G�%1 S�r��4��8&0&�"A)M{F�9��w�I��G��+�=c����.WX�q�_	6����O�5S�~�i�C2�]t�AT�.�_!S��T�k&����I��Ã7��ѥl����g������
�����0�"�!��*���O|Wh�*�x�y�*PX��,Q��s" ���[�E\��j���QX|n��i��v�G�O��,�����W����$�<��" pAi����`l�SG����5����wHkRI����OK}�(��b|���ӏE��M:��'f�1������aNK-�L3�e�����*��;44�{�7;�� *�%���Hc_{&��$Ϩ��T�U	�w��cv��|ʜݐ�d���p�%/i�[�!K���t-�l��/?�%M��Tuhn�?�1�B&BE�퇀.E�D��3
	�F��.<��<��s�	��b�X.z[����<�LK�Zm��%�%&��)��p��<����ې�}��A� ]��&�E
�:L��nZ4�vFB�Rn��b�W@��'�JX��6i�*$6����w�!ۛ��C�����ɀ����t�|�½2*�)�~��A+�&�#�'�'Q�dVcn!P������@��nO�� ���5��oZ�Ȓ�J��/ª3�S��֭g�֙���$3�֯G0j��{�?Te��ਁ�/%�|ˆ�'&���3�!� n|0rvz���3p������������*�;\OSٮW�#P�}Vc���Yuh��?�h.X����o�lVW6�W*pߞS��W�W�bl�]y}X���R
a�hS�6J;$��6ׅ�q�v����?x�o\�`ƵJ��O�#jRAﶔ96L]4\�/]Cv=�Y�c��+�LД��]��-*�lԟMd��M�ٞ%�i@���_����v����b��u5���Od�PTEd� �(�{�6�m��z�-1_���p�HpÛ���̽#����d��t� %b"@�`��*�ND�'SN�\I�t���Tay������m�S�����dT����tN�K6J&�Rj��[��������*s�3Wle�g��A����FcE�G/�s��<�A�fi��+.�S��!"H��`����.�Tt�[%�ƔMen�������[1���Vu�Gln���/~�?�&��Js�Y����|�4j�j��!�ؿ�4#	�&��V���sx��Ao�P���y��dX�p�a�eYoa��U �oo�Ԃ{~�$+GF� ��
lŢi��ʁ
�
���R
����U�{X[��;Z�S^M�_�t&b72�t6Ad�D���l�k�goK��iը4�x)� ܼ�������ޚ���VȽT��AO�qy�Ĉ59��1�-�F�&����=�����w�|�_{ht�����k���^*�g��Y��O��x�UA�|��c�V���S�:�[W�3Z̮��]��ږPNݡ��G�V$��}	8e��XIa]-���cbM���ǀh��ً ZJ��c ��݂&�JZ������1ܝM���2��B�m��0��qi����J�!8��d�z�&�fXb�}o���x�&�>Q�洖�L��}%��J
J8��������Ϙ��N���Ƣ�z�Ȃ��f��KS����E�g��i�Nh򼎹"��6K���}m=��Y�_ֶt���KQ��W��P��hsf��*�SRt��hH�8yT���zK��a�a;���4/�o��޹��'r.� t�Π2�;�S�:Om�L^�����L�c�QU���I��O�K�c1�B�7����L�9"���̛
3�� ��/$��3~�������薥��i���!Uk�<�0�M�Ȭ�{O�.��u�E*���d�J�����	��$*N�_5ヅظ���]|�t��1�XkU�}����Ъe��'�0���?�A�&�l:���^԰ j0�{���jyp�BV\����
F�^��^u���Xt��ב�d��u�p��]E�Z4iZ��$�g� �r���i���J�
$~Z�l�^�uJE��gc�����:�j�gkL�"���h�>#?Qw�>� ��z�
>����i���oMԏַ6�����Ȅ�'�E�]7�=��S�[+u�=��Uo���a��<�� ٕ���	<_�X�6$��!��X�T|��P �7�4��y�/&��&��>�h��JV�¨��u;�q�������`�㳡��^�oY���6������?��.�u��`����¤������0�O�[�z��G ���7x�d5�c�dȟ�}�Gd����u+]?�/Ҁ2�#ӈ	O|�����+�����2K��(�.�;)�r�\.�Fe�{��+� ����g��E�d�
�Gn����`}qy@^e=���c��N���<(1
�P��c�Y��A$�;������y�ㄬW�li{d&!3�%����rJ��8V��k9��/�xÝH��7w�o�SAzƑe�{���}�?u:Ȱ��R`�eZ~=rc����vf|��!V��@���Ƚ��CT[�,I�� ���.0�d{mg
�C��V����>r��3鳦�ijO�M�J�;�i%GB0�q��9���!�	u��?�f��SȿF����c�1��¥�M�!|zG�������^��t��_a�
��u��0��p�R۱�1B~�>�U��}��*�_�a���l��ܺd��w�hV6l�	ID+�C����:vI�H�熂&��_�}���X�rWzPF&���&�s%N�j�*K#���PU�czYtQfz�������iy" ���t l�{r׺@��������%p}�e�d.�C���n�(�A��:�-�I��s��:ѯ�'4���͛ٿBIV�q�md/�&S^�g���o{SY0�yr8vڇ�&�*�U��
��P��v��
j<�23��i.�� T^:���ߺ��i�Y��j�Z�0l]'����5M%R��e�z�?Ё��=/)?ܡ�@�}��v $�O�nT���_Y|��
�ߐ"�Ӳ���Ҧ7�S���F��k�����g�� ����&����8��s;��"�7�?d��-�I�~�`Xr�"�b5t`��ҫ���D�
󵼝���p�.h�whY��h�bUe��̣�\�����g ���~��g'`�Yg;X2s�\,O��|���v����X��-k����d���@��.�J��@{o�Ǫg����8��W�tEAY^�i"�n
�Q��l6�:#�-�8�K�y����3�w���0%;�o� }f�k  '�����β5$<rC���S�I:�p��P%��\e�)��u�V�KhB���N�@I[��"�/ؽE��G"��� �y����=0�G^�NP�}�zU���!��/�rҽ�qN-țP�E&��Y���{`�x��'�O'�F��+���j^����N���~�R)������z������.iR�+e}�+T���O6:?R$�S!�ߥ�}�_��Z��hVX���@��&^�c�ҿ�+�h}��><��.BG.�ا��&�g�J��名�R������(H��E��z�)�����'JTs��1��'�L����5�,���m��ϩ��4�'M�C�bY#\t��P��:�2�-H�:�T������+�A��*�����|�pKL^,��u��6��+=��:!���ذ?���������+t	q�:�78;Y���¶p24T�f�}Bie9�uwT�b31�a�����\��Am�_R�F�3���p��&�$��h�!�����V&��������D��p2����ԣ�����p��>C�C�Z�!H?i����ζ�����T��Vs��}�Pj�����iρ>u�k|X�i�20���O�,�/�jNXu�O�g��%�?xq�iڻ�ȼQ�>�WN�[J�,a��oy�P���7߫m�E��s#䡿��ME�VnA�Ý0d�{�
OOc!G��� |l��@��lˌ��k+p�ۥh�L�Wku����]c�x��̫ �������g���i�|I5�h|?����H�6�]nI�1��U���YB���:J"��8��< ���q��/�������H��$�'?��t��D�	PB��CM<Wt�*l�mg���r2<cFu�:M�c9��闝ۑC7+ݞ(���|�Kh5�u]���a2i!���e�C��|x����rU�b�7��XL�r\����"?Kċ"u6��E~��w��|3?a��H�4��}u~SР��lӺ؞r�=�Z�a��+N�X��%A#�b\?b�����H��@<�������h�L�k?�Y��z,�i��9l�(��_��A�g�C�֛�5���9���u��\��R���w ,�9�w�a���E<vΈ���@7��z�Qa��{0ʚ.(j��B-$%u���1˵W�濋<ԟǏ>	n�YeV�:;���͒R��6��F�g��� ��1�}_�{4��26��OB��ez�h�dK� ��PH�n����4M5E�̨˳�5j5�b�w��n����L#<�d�xtLl�����u10,�[�;c����x��%�$1ҝ"��%�^4 z���ĖY��Y�~���=��h�3�'���eHϿ�e�1:"y%- �!YF��@T��p�Z�Z�ru�D�A7�1"mfz��$��1�]��^���(<��W;e�;Ϡh��9��E3� !���,�$����{88���ė��qj�#���Z���<[s�n8�Z��#'kp�1h
�)�q��N	ٛ����nu�T�R: ��?���2wŽ���]�����i|��2�;�����[��W�m����_9��M ��y�)$�_�c��2i��B�﷬]��d���)R�Bv��V["�8�^_��u�6,<��46~⑀`���I;��s+N��/ m�jՂz��Em�Ɠ9ީ�ڞ^��n�y���E�&�-�9��& ^����v_�\ß�xzd��t!>6�t�A��'�����r̫b�8�jm�����E.��u+q�`#ܳ�I�]<�\ʨ2��* ��e�ɆSߡs@%U��-*�?{v���H��_���[�~�9 (���%�l���S�$�!�z����u���P�"R-'�ݽiCT��2_�C\��!�Dx=�E�\��y���F��-�_�0J �HbZs��*F����q����yڬT
�0d��Y�#��\V���EA�_6��EkY��r�����u�O����a�,g�Ș~Y)���V|S>��x�����R���Y<l��������W̥[�̾�~;�u���Zd?/�� :�m��]�9g��4�藳���5m�O�'p;$����b�+�s���>�ϊ�T#��冷�]5_UG�.��՟�zD����9��hzR�v����\:V!~lӻ�a5H�NO������2+�����"��.�-?g��z�:Y�����V��h�l{!�E�.�PR���vIVHQ��*ǻ zo�*�V7˽�SF_m+z�d�O���/?���g�0c�ӰT�O/8X���[(2���q�a�)�l������	L�S��ؓ�{cmJ�D���A�qkD�$����%���$C0�b&�[J��q+:󫬻q�9r����9��>�C���i��7�l�qU�3���3!��Q�tJ��!�Φ"�-,�,��t�X�2ѥ�o�v�5A�׈��n���� R��H@+�9����4G6ˇ���`�d��R��]���%S��C��Z���F��tѿ$ �+��f�
���,�z�]Ra��HE�� f-��j��'���I9�PF|��'k)NW�D�6�iV5��Y�4_G��ɝ*��Xɔ��a�C��|����A�jBzfy7�Ld�������T����m�B+�D���8:S�\���e�8v�|�5����FH������s�3j�;]�/S�ո�sKu�������O�h�W6�ںu��+ֱz�3\ˈn0jSu��BӠ�wI�O�*�Y��.x�X�s���Zp~��[z?�#nHQ���0љ���]��}Ň�`����z�,���˽�H�4���"����Fͨ���P�lA6�9�m����O�?�����1����D��}����.~��FԔ���fĒx"	-�������B�y�큎H� w��I�zE��h��v(���0/^IE=�&7�$������8�H'w=<NF�0
6@�5S����T��X̣Z��U�	ӉV�y�Uy"n�է2���G^��P��D��jl���3�oe��"��B�]�,��:B�I��F�q�ʩN�}��.�^�/�O�!h�kf���93�A�>%e�J�cP�4K;\���M������8;zX�_;k��h��.�(�4#c�a�Z���)4Og��̬�Y��P �y�I���������ڠu��K!����	�_���ݸaf�W��9�^^��9�'X�^��V��4r��cG�
 �e�Mni�"�d��J�~{��k�����s����`��>O��mn��㸬��7�T���w-W���&D��� ��P9c�����@��<%�u�����e'�FטF�0qH�R��/�D�j�y�4�}��3�f��i
t�D�2�a�(�� ��/�(������J����p��Ğ����8��9��c��j
��~fl�q]M�"�oKQkB��"ѥ�p�7˄4�'Y|�P�9�>9�hOc/R�?����I���5�s�������F������$֫���{6�3Y����.�Q�/���o�h�3�;O��Y1�2�c%�Y�N"�3�82��>�{�W��W9��Xw�1�D�s1l�J����5+c���\:`Ϛ��%��aFZ7�0z�'Q�;�
�@S��NUD��q��p�3L��#��-/�\��_�0/q�5G�/����B]<�DSowxݻ"��+l�e2m�ғ���v��C4ΒMT���3~�pP�p����M��0.���O�;K;���B�<zE��F�oM�߮N�b$yj��'���풋�(Rn�޼֐�P$}��	�������+��M���槳�[�̶��b�]�h(-!��`���b^ȉ�h��c����_d!8p�Y��9��'���*������F�AOP������_0m*�[���3T�<'D��̃X�8kΗM��vI�j=�9�&�i+;P�n����A0I>|ѝ�g_d��x����?�ߎ�Q��`꺾'�4��AsJ!���
�����DXX*)���pK��>|�KP�
I����Z�~l�^�Ȕٗ�c�TYR��$輨Gx/K?�A�\�e�Bl��d伟q"Y���`�c|���;�o��\���x�N�I����q��,��~BK:Q1� ��K�8�3�ی�oZ��	�G��:�z?�����	�v#9� k*j��73�c��tKm�#K,�7�����D���d�K}��i��|ǀΊ�T�5�X��N����*e�U��M:iٗ�y�(Z6i��P��|d1���������!d|�>1����gG�y�= Ho=��ԘK:iK��{y}�t?�g.��
���+�����_�(`kP�AϙIR `<��~|��K��;��m��osv�JN'Ǖ	�V�/��'�؆��re�C����oL�BBb�{���O�'Z�*���P��ڶ�����N���X���|���مp�#�	��\��[L#B��a=��C|C�S%+�eΞА�v��Q�6f����G�C?�͌��x;�H��A	xXo�x`4 �n±���S� ԥ>���j��u��y\m��j��I�&���㇙�7^uu��0�P��W��rY?���0"1��q\UJ)�rAt���c'�+ڧ�jR��n+@�c���j$a��C����������w�I��\�Q��]ڕ�Ǯ����~���ruU�YOO�#�����!����;���q9��g��`g����[��n��9��|b_ۊ�,aCڲ�iV��_��/�� b"�m�%G���?��.o�7S��<���]��˰�$[B��Gk<|�y�������/�O�s%Yb��K��4�cNو,S!�����P^N!�*��g�i�W=�3���g��"q�O�M~������@���<�����o�����	"6�0�����@[MF1I����]����Q=�KN���=���l�����@y�YSek�u�^�2`7�+�������N�h5��rt�a�|+������o�X.��0Q�"熀6�9�T�/Z��(x!��lEM�2���J�Zp��YE�ع�����P+��t?�]=�P�b�dII�����1�E��&a�'jCґ?^�n�b0������G͈`M+KF�3�ի�_F;u;�d8N���v���vJ���Hl"pl>��j�A��ԥ�o�ZyeI�>�?{d��d���ǔ̣���F9�K!��s��n�R�d�J�Al
�� :Ֆ�㭒E�zz�4f#�rcݫ&\$�[Eκi�X0L;:m~#��C|����o��G����S@()���p�&�a8��\��R)m/��"%�\�A�V�>
wQrV�}H��/��S5��C�H���R2ӕ��跣a��'>���hq0y| �8�����F�HWX7m�������$ob�˛Z��@��X�XK����24�z���,���kQ���Jah��Z��^t�jb�0�<z"��](-�w^�����YJ��T��72��-���Kb8W���թ���S S�;@o���t����<=���{��	D{����	6��c�_ed�b�oI�� P�vs�rQs��w*�A�� ,�p�%���>���Yq[�g?�f#�S}�ǐ&������ޙn��ھ�����.JrǑb��ѿ��0N�#AhMv_AOyFt^�E�Z #0t����ޏz�~�;G_������a02�N^�'<�=�)�h~���#�L�G�Ս��~7h_�⑩]d�1��Ry$)��Q��ə%�.lP���d���
{�a��~�ɵ)����,�j�`�O2��Jʓ�D�m�[����^' 3+ĭ�����-)�I-�{ ��O�[:��C ��7�&IN�p�x�� +�w)��5](oϮ�X`��y6����"
|���#���@�� ��**����6e�z/О�CsΨ~����,ْ
˦	+��W2��%a`��C/�2D��Q-�b6��U���[Q0޿I_���[�X�O|���r�I،�vi�|@_A�r�P��U��aiY�?v2�;*�Q"I(*�G����<v�Z�@Ga^��F&�Y�w�jToi��O�̏m�(^!�&�g�_��}[\`�.+�6��q	v�=nG-=�P,(X�S��F�:oWt�UTHu����&���P�C;138��;�w@zĪBl<��eѴn75O���N�g]�%��Ƒ8pp#ݓ��\�~�_Ly�?_�҆%ӎ~���1�I��?�qU�#E��f���f�+@�҉���B
tM��D��~>��:�YX��.�HGU�L���Z�I��7NH����dKci
���+��;�{���y�![���J� f�Чl<a��m'�Z$
`�~�mj����Bp�b�櫲#s�Q�>�tDe��`�Y��.E�"el�s!���$Q���w������۱ˁ�ɋ�ۤ	�7CKZ�rA�	�6���Xe�l{ ��Pը�$R��J~c�\:"�t�yh��J\߁�&(a$����&����� ��#�|A��m�O���_���;}�}%4 �7(�X�[�9u��!�&��g�� �
Rr��1�F Y��I�27xH��ZޣP-���� �T[�G&�=��ݿ��y�yU��r����Ґزğ�.�xiY��j��Y��)�qDh�9:%� o�����������p��6���������v�'jl ��<~+��=���M뭟�sC�=��9��Q�"t�d~!
�������-ۮ�Y�T5���b{EN7Gs�����>v��Zq�|*_͊C{�F�~��)��N��*?G/��+�X����䵞"�S<[��S�ׇ[��+zA�Pn�LrA(��l2o-t:�I� ��" �N��2@ߢ�_{�hB߼�x��Ԓ��EfJ�0��=��"�b��2<�7A����S��+���X��jL�܋�tC��VNdӌ�iK����cI�����]���'�Pyf���+u˸���t�P{�q�	$,}G������L�I�TR.�ZQ%�;*=-\��s.�]e��:N�U_ѷ!1E�?���sW�!�Á8�qLn�,T����=È�B���`�O��o�S��f���I	#4Z5H�[��'#_nl�������O�����&���'r���`^�̴uH,G��(w�\��{�ĩ�cF�r����$!&�K�K�M��l!4�A�K��S�+.%�
|�ʥ�+��b�7��ߊ���[�r�[Q9B%����ⷢ���K����v��l�Q^Xk<��|啽����*�W:��,8��%Ҥ���!�1:-��2���Y<E.�C�F�VՐ�Zn�a�n�Av$tAv�v�'lB�&��7e�i=�&����o���3��~�j�9��q�[2iQl����d��s�G��P��3qSP�n�A@��\�Dw������_˗�/[�\�S��	�`r?:N,M7:�B8�q ǃ���S1�B�^t�X�!��R���\��`"2��ة���H��!A�X��	�+����O��:����j�����P�n�~GgX���LBy����'�,D;}:�3]=��Env6�Ud�g��pa����]\�-*#�$LN$}���5nF��8_*��Hh-��%:?����-���RR�1P|nZ� �;���b1��J�D;aBzpG�V�G�6%T���Bs᫗^�<ɛC�,�,�54(��i]�����w[�Cjw����B�h��x�05��r6�Y�Y�Q��
$ڪ���$����$B��E}h<*_5d	�̖�8���k�(1{y��̰�A���C�,5P��PE����"��J_V6.�45����P.`�]�é���Y}�`D��6Du�m��Y�0���F/�d��dJ�'�w)n�`6��N�Ǝ):(����� Jp��+��*����4�b�@lO�$a�S��z��h4wj����z �pjY�RG�%Xbx����1��(���s�߯p n�S\�n�b���\샄#4���_y���C~8%�(��b+:�K�h �9z�$�M^�[?U�~﹅�t� LF��((��}�Y}��Ջ��O��@����~~�=
S��o�I(��o�������7싈YB���h4��z��8��y�|
�CD�*�ʆ�B#%2l�o�f~!�%^�}U�����a����q�I<@E@�.���9��#��<�8� ��nZ-!����F���&��-�l�%����{7�e.�D��q�lp��qٹ�C��	y��r���a_�ٔ|� -0)����nMdOB����5l����3�8ӿR[[����3pߓl��Ч(|x/�r��c$��'��q�P�X"���R�`���)wl�n���r�i�Z��E0=�/qm�J�`�)����7z!�ye/�'@q%s�k�@�􁹢[��%���oYڿ�g�Ӗq��7�����nZJ�`�o:򼳸��N�������{�%T����_&���r.��p�h�#�ٔ�?1���ӣ��%�ʂ��6�]a�+�6�8\#^q��~g؂���@8��8B.c'n��Y�=>��*q�?��~�*�ޤ�.�i&"���X�T����Ɩ��:�|�����za/�$�S[���R�=�x�^G�n6��4�*����s誕��(9���ۍ�2pݕ�M���}��荨[�D��Ɨ��t��í�2��G��7�����א�6A*�c��\h����NN:���,r ��COS������q�)Qq�N��C�Y�������:�A
"78]�Y���(#���=�!� ��}k%��9I�Z$ 	�h�?���m��@�U�
�%y�odzu�'��9��KY��ɑg�1������N����C��1.?2k��"{��9�6"�5�ӹmO������������g���Y���S��lf1��	�n�����k���&1ұc1x��H_�$<@M:��E�r`��X7��z������l�>�( ���R��K##�.�)_L�����D��\K���Ȉ��ev�G�١�}y�A��\�U!��Ρ���u�@(�-��	�h/�yN̰��>�1O���������o�^�"��b�A$̡���?�= ��"��`�����9ΞZ���էX����#�1j�0u#oC O���`m�d���m���%��%�A�%c�6O��s�����H�s�l��q�>��A�B��W�yj�!HA��Ŵ��2��D�W�5�V=i���}L/:�T]רV1�|�0t�xLԠYn�:^o�k�3hJ��gkKnr3`���P��r�l��50����ĳ�Hǽv&���ފ���-M_I�pM��|��A��`�7��y�|N.eH�n���Xn��������f4Zt~r�Gn��F@辆���B�@�Eu!<�vi��嘛LBm8ï�{;����[$��J%�}�>�������U7\Y���Z	_ս�F厺XS��b�T+z5
	%$̺Γ�%c5q6�)��V8o�ߗ�\�t��!E=��S3�6��ɱ��-,��̔:-����_C/��<��Z~'��R
�>�q[�O�P	Ѱ�|S�j��!�Ԫ����&|�R�	����|Y���d�]�2��C�<x报�c5C��1S��Cw���GB�T��� f��A�T��P��T�<�Xl3;����5�*;D'��]�\ƺmUJ�:[��?��(x+��� 7Z�t}U�-��s[G���%/r��k(Y��8M�M���?�]q��y��r�B�A�0�fȗ�9c�Y�HG��7���oW����/KaF� sa)�+׈8ATI��CE�������F��Ơ=uRSI��3�����w���H)L�Lc���Wx�
l�?S5�W��@q�!6ί�6� ^jL�>h�5L�E��>���2I_���B�9�I�ۥ��������>�a[#�����?n�(��WA��tY�g��p��� ��/�5u pa��@.E���:�����&���3�Q��\=}�aMw(*�h�oD
�*+�H�� �#�lD"��ʕ���w��S[[�.�&R^�X�����Z���-[����Qv� �Q�eEң��e�֫��u?Ti���c�P��&T�������`gyN���B�G��?_������l��Δ��������ֲ �Κ/~1!}/���aGF�w>ՀA�B�\�П��S!��)c�߫��Û;�HX�_O�E#m�M�I�Ess������;�m�?+mKJA��ͫC��κ(_T6�E�Y����t�O�A:����N��%���Q�г 6o5و�ڇ*~c��H���Y�۹�d�m)މ��\"��D��M�X~ﰦǳ��o;��'�KH�Ι��R͊�Xa���R���ah|{J2ϳ��'t��ݡ��ɵ����e��>�,;AD0�U5�6��i	K�t3���}k5k y���A���v,����v��MD,]�6=7aԬ����`��sY$;��FR���c]ҥm;5Y�P+oA6�T�oh�Lo;_�pu!RO��3�� `�����A'�گ����w��2���loH�0�82�!��gG��}�����%�Lbn�E�����MX:�j����z�*,������N<.&%]�x*���J��k�i}[���j?i.B�j��7�d�Kp[eHױ �PM �_ɰ���+H��,;��b�*�7�Օ��H��Z��$�ԕT�ɶ���6�J�T�4�}u�&5�`��8�g����yIo��B`�������&����k�w��]N��'R�_�WU��Zq���Z_�=^"ќ���#� Jgyz���9�r�cd^�u��ə����t�4�\.T�� CM�����y�0݌r�}�h�YȢ�cH�B˸���!e�VD�>*��cMV�_����C�7�QbqU�(�Kh:�tS<m݌N��Bo��(�Ä�N�����LM��y��2�J�F?Gܧ}���Qse�%V1r�x���Ny8%:��eY��j���]���������)����z�]� A��Y��iW}��ݐ3�B�&�ۥf����@ƫ�&����e�f�<�d1e�W�0�I�$�:LZOwX�?0d,Pc4u��4��u*�gQ�v�z��`�����4�)��!dR��&�%�H��qB?
O��P>i�P��_rz�H0\�1̠�р����`^�N~�����X��Q�b�G��s�
R�K4[��Qя({*�ρ�/6�����nIŝH�M��-�K�B@d>�	�
�]F�i��i)c����~�|��4L��'�+֖0u�E��gƨ���?���e����:�n����NPM�W�A�N�xqVn�	s<�&;�1���f=%����Y��W��J.�c*���X�I����<i�����k����GSôH~V&?�ܦ
����ب�"��;�	g&�&b��`�B��e�c��;�l9_j�����2�r?�����@ʷ���S>�brQ���9�]���Y��{�`Q�_=l�s�_x8�4�!����ҏ9��"RaJ��Y�GY�,E�B��O�z4&�Z25�����?v�� T��҇-�.צ�xSh7)�)�	S���Z\M��~r��*���b%�b.Ƃ�|��!�`�z�J��nl�{�A8�I!*�����Sa��9A�+��1�H/��?9hQ�~i�B��<'h@�L&f��� �6�\����2p��ǥ��-�����8=��I����	!�I�$p�&gF��co�ګ,T��:f���Q�A!�~@�R��?jE���.�ض�<�A�|��ـ8Jу>j�3�-��eHS�Z	��-����;���^r�=:g�J�#��iǹ���:��P!/�m���䞕@�����lx���o��E�f&'�QW4�[}x,:!͏�W�^��BPŅ(:��A�c�y9��[� m�S.����w��˵}�dBuܗJ:�H\ę�ky���7<�(�:��)���]�lۼ��x>�D8��'#��خxߠ{�R��j�1k��z��0�)�%q]�.g�̏��qF9,X���(x-��NZ�Q�Si�s��܏�w���%�Ұ�3��G�����0#���YC��#���&K�5�7žq',�,���@**a��c���QC ���'|�;s�ޅr��;S��3i"0z�N�X߸��[9'�\���vz:�8xz�^N`�)�MՈ�'|,P"#��g�D�{�����^�&dc� �p+	,E<�J�w���nTt)��`�X�
$�K�X|�-�Qv������w/M�K��r�(���1���Uo�?|��_��/��|��Ҩ��ڹ���{&���x�;v��B�
��RpwJ��k	�Lj����Ņn�'�u��n�|��s%O�qW���~�����$��p�֔�C�F?$��u<ؐ�R::Nz��G��5�鎥`���)
߂��S�O
ho��=�K`B�_�3�C��+�����iK�{�*�p��M ��V�1 ])��X���m�m��I��p���i:�_���W��Y�mǥ�R����*:i�mG
[! �dMw.-�q��x,����GM�����s�vϽ��[L. ��r�KVf���WAE��W�H5Aw�`�=�����f%h޼�
`�y�~���κ��AB��⅀�':N~]�� ����`?��7($��8R�ϱ>�,`�oDـf��3��Gg���S�o���?iM������i�����g�#��@�>�k:s�nX��6L��*59O���m-v( ���)�Z%�-u�4��r�u�
 ��f'n���������/DF� }�M�t��ƿO���ت�-D��1 1�u�����K��e��X��,7�����e��◩)~��A;R����K���Rv#*Pw��5��U����ԉ3V����uR��y�ǎo�A�-�O$���N������$lr�c�V1�e�t���Q�/��zj����r*T6Ie����-ga���+�[��#>m��ԧ����S8��a7$VjÁbF���q	��KF\x!C��/yb�Vtܓ���	� ��_�h-���N��t¼���i��RX���,s�+�z(�g��y�"1_�,�"�ԉ&���%��A��:����9�upt�����COWH��u�l�DϟQ�T��$N:���Kу_��t�_S�1й_�}��nTGwJpĔZX��=�����:/���	�����%Vx�4ڵ)���2&��q�����vD,�>1���^_���9k f��~/�W�zHf���������`X�R;��7�)5�+'!W`=P#�M~ɴ���M+K>�A'�	��J��+��%i-���1�g6#%t�v���(�'�S��#A�Oi�_OorD������&��1'@����0���4QA�F�0��?���QI��MY�wr6��ktbd�g�>���lk��Dӆ�U����$��ҍ�h|=DK�S|�&%b��@Z��0��^���<��M���h,l��rKŭ���:��R���m��h�KP�e�"�ЖcNY�"ce��/a�F�Z�t5�J�]�&��R�u
ir&�w-@�;�ƷjDD�Cj�i��A�����t�|nQԶ
�Ob�n��=����$�/ı<)��)�:�+����BȨ���<�����V"r�®�'*|��V:�S#�8����f�(-F;3���|yZy���)���sv��H���ķ�U78����9�����N"�����Q�ez$>d�5n^^K4��t�ۥK�;q����V���9E�Ɠ7f9;�������0�z�v�p�N��Z$��-�x,a���s���W`�O��J�`��R����b��O��p�<
k.;_	���:~�g�/0Ͻ@q��y�@�!,v}zcY�Z��5������<��:�[˱���4V؏���Z���%�Go��'.g�;�mX2\_�`O���i5醼��멑'�v������:��	�k
��)S��e���-�g��M�2U蓀!{�Y	�?�w�U��3|�t�*ȏ̷�i��T���|U�hm�����ؒe�+���d���^�Я�����jZ']�����n$�|�M?Q!�}Ew&EK�������|L[�]��!��2&%��N ��?ڇ;�y���G8t�Ϙ9��G�L�8(H���4nQ��>U�<����=�-U���I`H����#�mK�[�bi
(q�h�r,OT�P�����twW����P� �p���y�~!("�g�)�K����%��1�̑�Z2�-W.���T݄8N���L:� ��Fb�֢���&pB��9�����;�����vM�7��>�S�Y@���� ����-�"垫��C�V��
/�.J��ʼ9�g Z��F�=Fg���
!/�`%#J��Z�UW),Y8d�N��N��WVݬt��d<�Z�NX)��4%@�9��!�Z��;���j�?~(��g��`�L1��E�	���-�^�>���=���Tى�Nb4�-^��!ϊd�]G�X�@$4�1W��STJalNf,�����I�,�mȸ:ҷR��eG�i�c���,��A%i��*��L�!�Á��@4F�wz��scZ����U�h�喰p� �\'IQ�:��H��[�=��4?���Wx���:�Z`4PS��f7�]���KP� �|�=�T�j�m��#<�ӑ8P�~�p	B������Q��r��5&��.��
��tBf��!��a�(�95gx
�k�K�a�����$�6��}	�c�j��״DZ^M�~$�",�7����Cz�۟�(����}3	{��эut;�@�诈���l�ޛ��n5v�]A�~.�B�Yn��U�&���䥣l�˝��BQ�4d�YF���/�X����t�=�h�uN�A���)I(44�ǒ�67t��"o��paf��|�w&w��06R.Ob��l���Sx�>���7�y*z<W��d)zGG�E����a3E^��U�7e�~m?e�V�2�.� P��,7�_jI�0*L�g�ƃ7�K���P�﬜FS���{`ڄ�=W�O���q�M���!0��[�H�f/��Lx�J��B��	�0�GxVK��K���<�<:�6e�ivy��XW�*��-�\�V�y���*0�viжl0T���m����<d�I|$�Me���1�~$�}�p�Dݝ�`	^��d��QIL���NTO�;K*�Q�#�rgoz�K�+��_\��L�������z�k�Ь=1��FA����<�(T'F���9j���H�Rf���H�H��p�S�"��|2����|�ZO�M�LG��g4;-��m�WV{B�w��we�FHÿ_�]r�s4W�C�8\vR1���������#�N�8Y`���`�&��s�T��`�֥����L�X�&Љ�W�"ȩT����!X�(K4+*�})�süO�4t^� �_�倸���>�BF82�5�v?�n�,i	v���r�91�7"LAb"��`CU�kmyDƆ\) ya�⦌������P%%5_LXGV��HL(6��vA+
#�AUt.0<i&�?��ln����,yY�����؞������u�(�1kd ^�s#�!< N��J}<H 7�f��Rx�MK�����'}�����&��YQkC�)^E��;Xe�[>qUF?�-H<&ڝ�?��&�L/����ё*���}[��E��T�i��N��3⟤��Gz�4��EHn/!]I�k0xy�l
#Ŗ�A�|�=a��[��g�q��se��\ҷ]��5����L��z�^�ᕚf8��������]�mv:W�|!�WC �jr��+ �@��dlx��7B����Mפ��k�1To���������lOz�4��6c;��,g�����څ�ϋ�
Oؐ�M�$�(Y�z�a-�G]1�f�}|�uJ݅��n��c�a"�{Z���i��ڇSL��Q�P�3,uc����T�G�VJoP斱��Pf���C�:�κ��3D!��� �4ͨ����	#J��)_���ɤ��z�f���|�2���E��X��,����z�3(�0)m	f"���w�D��b����y���2+-Y��1f�88���e�~P��E�@Zg�*�K�.u�,Y�7g�-�W��F8��を�(���3@�Qe���υ�\`�F
��{y��Df��*T��h������AJ��������i-���{m��8?^k�`@z��|��5��;���fs���kv�.q�ro���-UZTg�iS_|�iP4�| ¢qL����������;2;��Q���Se�\L6N�"K4�Ş0��=\嫦���Z�/�q���ZZ�}逽����׼�N^5��1�x�	x�����woRe��dW��	�(�m���7�L�_�L���)4Ӡ�㾼��,�͈��2Ҵ�A�����||�}�f�CZa͏��c��1�V��{��i+���@3��Ħ��[����c���n� b/�gW�y�-$���A�2�{���R'�Gb0H��[^P��B?_��ĳ��y����'>n-'�7Q<�1�C��2{� ���Lyd�ħ+���.�y��귡	��AoW�k����l��-x���-�a53$t�;Y�b1��"�hA�r}�����YL:߮ujj�hXT���31-B���ε���[1{O�{Ւy��k��Ssk��}x����}Gb��u���hOԆ��Ӯ����h����K�ZA}����#��b%�����0��o"b!�ѕR�3�g�nOE�/�N�д��Z�Pg���U�%.��5�{bF���G�21�����ka�p�s��"֘�=r���_��.%EG��Y�P�]�.̜���+<�m��9�;)�_���CF*%�k
��<*����Å`?�M�E�8%�v�0K��0���P=������A��X:<u�>��_$9���s/83��ﲯ\�s�M;�����b�b�{KF%|�*�%���׍8u�[���0:f$er7D�~��n�f�X�"�p��5��!�*Q��M�߱6��X9u@�`�FZ�%*���/��D��
�����%�����cj�5r���'Z���92������?5���l�k`����ر����T�GG��j����W�;7��t�>r�O�)�|_/A6�cQ�W+����K�rrY��:O��(��B=�L��n��igS5�H��x�s�ɋ�*�c��*q�_��N*J����gn@o쐁Ki/5�ì�u�٪��|Bm�$d��wɡ�̷�ީ1�/K|�pKr|������?�ky5 <n���N Nguf����u���m8D�cp���ws�fy�p�ׂ�(|��ζJȕ��Q�,��96�qz2���c�/�KmW?��v������FB�&WP�r����?chׯgҼ�6|J��B��e���(�>!0�Ek��M7�	�\Z�`�c*�`�Q?֌WGSB�%�"0{�drI�܅����rU}b���ͦ�ޕx}��H#��_3K|窻qD=��mi+�Ё<A���cM���D4��3g�Y�r���s�%G�>Zd_)Sn3�ޡ��{l?B�����c�����-�Rs��2g�����8�[T�ۣ�^�:@��d����b�B�&��W�?;�E8Y H�eͻ_���4�?�����bV����=�[1���Q�l��-��.4eM1�g��1�D2�8��T�vg[]�@���m�WY�gM�y��!��:�94�=	'T���d"�FH��T�ӫ�UX\��Hw�"�82��Q���m�Ooix�t�Lk๮k(��{lEz�<�Ji��	��6L��ş_�J�WJn��5�cxG�nw�N����Z������w��%=@��H�ʇ3/�� �t(׳�z[�܄������eo�ݛļff�D ��U�_��&�lޮ/`��?�p��O,N���g؝�ƿ~'������ �@�E��8��1hE?������k�<bi%tʷnn{���­��Ly#���Vйd��s��)��Fy���8nZl�!�s�<������V�=ۧ�ԫ�+W��g`n0��vw}����N�JS3��=f�܄�,h����sd��~��d�W�B��j �؈����5��I�|�[I%�.~��" ���=:�}Q�������9�6)�&��/��"����x�3Gے�[V[95��r"�D��F������,Q:��|p�٥����F?�f����>а��w��LU
��u�A $Xii�=�`��Ph�ʛ�Ty]��b3��A|������G~�>/N� �1����"-J�ˬ��L~�eK-�&Oժ�0J�#�����~�'�lb�UcF�����0��}=�E��!?���|�?����X�!���^�<��YѻMO�BY4k�׳ Z�Mѧ��T������ZP=��U���#ڟ8ˆd��nL-��~/�G#:�n|������T�;��JJO^��܋Amxo	:imP��.3�7�MJ�ŷE�v�?B/~��FJ�R��1�6P�8u���l!�>�\�@'!a��6�(xX�]��Ҩ&�O�l[�K��[�P59�L�L�
Bfho�i�HS�dV s3&9s�P4]"�����5}z�`�7�]ŵ�^vd5ŭB�{$?���z�U�N�.�|����#�`�6Г��֢����i�L->Q2S��2kw���O������	l1^���*��������@�w���Bv��a�JC�yE�HR���2@��� K���O�ac%����锥'����-�j�0�p�=�BXox�^~Y�!��J
���ą�]��C�:+�z�
�0LH��X����:�g!�r�d����َ������rNL����d���l�?e��K��_b�RE q��V���ߧF!�|^2w`����r���DĒG��a��G#�[�Є9x���q�6�ci�/m5���T���PG绱�{COV�=��,��#;yL��N!��R��*��|5x����f��LDLq|םzw��,��}��wty�3a�>!����G0��Bƒ�L��g���B�Db��cQW޿����4�?���T2�`Z�����9�&v��a+y��/�m�NÓ�f���m�@K���F�WԖ���2�`�OH'7�JktR'�`f�*���
V+,N�DK��x�����%O
H�	�/�W�=U(&=�P���˰������7���*�:�7zu�����	8�|H0cT�9$ᖌ	����K4'��=�+���lQr���� c�q/<>�s�b��S���%�N9���ul����=�>/~}�ɇ�բs�H%�*a=��eY��֣�wCw���8Q��W�,^�2�L�U��?Pa۝XK	�k��u}��$����O����t��6��0�z�a���hg�2�6H$41���`��?��u���̓�m���ׅ?�x�nXB���Ä=EK�2��m� �Ti��-?�e��{�F�X�5�ax��+栫O����&Lф�OV/����+�W^��d ������03L{��Vi�Z������2�N��ؘ�q��,��K������T�P�lDW�}�r@���aq���²>�_�iw��IL`	u���v��[�DN��lU�d(P�w�~���,+�M|�e�U�� ��m~?Q��L8���}��Z������u濽�z�dךN�$ﻈa��&;:��ýF��.DN����Z��W�pV%�����}�b;�#g�!b*l�zY��^��պ���u�bQ�����դ�Mc���K&M��| ��%����b��(�}��/�LI]Fg��]�\l6�0�����T8���0E6rq������U���+�,S=~-^hI�F�x��aƶ`�^��d�?��n��q��XQ�ͥ<���.m�� ��Oe�#����#�x<C:��R2]'��*0�f��	�Ʊ7�Xe��l
p
��1(�y����K�������ՠ�-�9D\kO�v�����t0��uҌ����̠=�!��Z�su*��Y@��{D���'�6�n*&_�L�xg��qV4�7����
���iz%��d:	�i�`Z��l4ׯ	x���_�.12k��u��y4}�p�>�I�`j���^e�%�҉}9�:ʎ�p�c[?L��(��ǉ���[ÌC�ZPQrμN����U��8��n��!NK�
�~�cJ[m}�.[���gJ�Y��|7��}=䦦5����I�O�u� �r���a���pX�]/�J@�>�q�h"��.��|��YTu^�i�-��TL�~���� ���GX5^4��Lz��+�k��	h��C�~޸���HiK P�n���	=Ѯ��;��� ��/�à05�P��cTq���d{�Gfyg�3�%Zx�C�y,�'n�ݒ�K��е�r��{�rR��&���sCV���Uhz��hHp K,�#?6����}�%�r\x@�1�;�;e�0���=>�/��X�	!���7�bo
8�9�2�H#�x��7�F���91�Y��rm�?V,���:�;��{k\�,�������vOF�U6㞣�����7�Ps|�u�L����s0�&`Q���s��c��=7������[6���"up�@�ɳ*I>�86����pA��s��X�E]$��֤`3U�_i&4/��Ϲ�i�uL�U�c�G��+�LI�"����^[���O�v�`FRg��c�Y@�-]������#�(~��gy�2�c�W�ߌ��W�k���#omK�̱�J�Oɺ�n�:������+���l�<1RChg�.
�7�#|;�A���}�ʨx;�dIx�Հ��k��u��gf����NHHϜY��fʻ���BG!�f�F]���f$���ᕤx����Uւt����7��"h��R@_�6aa�;���>.M�E�%�9��"�jT7S�n_�r��g�\�XMv�ŗ
JdGL_�h� �)l�l.f��6	�6��5�=��[|�#��}�8�	��?K��c�N�����~DU��_�Vθt�Qj�x?><6��4�\��[�X��:Gք�y�'�;ۜ~\���?rq_���ݭ.�#��b�v�Z�E��� �Ȼ��E5�k����l�s���h��)�d:>���y8����t��2���h]�<��_��F�-x�6G�CWt�.f0!e-�q]]�'�!���g_Q8(=<�Ov.�|�RIʦk�v��	�RUG������?-,Y���[S���Yg�?xa
t_űd�q��Yֺtmm0@�ǑK��{Zdu�U�jA�q�AO^z-����e�� ���D�w�|��{͓M��(N��̟�U܍-�A��˒ɵ�Ĥ?[��>Ag^K

l����f�oD��^�;��5�I_YX�����~ Zp����;Tf��?3��"Ү�e+L��2p�6CۑXH֔�'��3趆��m���?���U��K��(�h�h|��|��:��)�`�r�%m���RB�˘�ucxU��4H�"Y��a�W����&84��2\���t�����#�SX=��l�<<ڪ�0a��K~��e�U��lE5�l���1�ݧY�^W���[�*�"Sn|'����$H��ğ�_ˑQ�i6��X��%�@���,��/����6��_6�{R �	�
r�Ө;�K���'��b�	�Y/�C�VjDF6:g�}"��}�6���3��3k������J���.�
�]�3t�|�4^�f�H��=zx[iF}Uŋ��gC,���nt0��wf>W��}pz�'����YU�m��誐�.*24�0Y�5'E��sU��un���i�w���V	o��&�Wo��U��M}X14���Ba���oު�#��ZҲ�V �7FV��ɲ���?��:���C&�,2�@������ܑ��>��?�:dz![D�x|���
B��)],K������J=/�F���v��^D�s�8��j3e#5��X^�6��:�VͮS?���?��MY��s��B |MS� �@�o�
i�C�2�LF
�"د�:�ŪpQ�/�'ν�wS�%�-]���׫�j�oN�ZӢ}H�m�ĕS�٠\�DL5ל���ܢZ���&�G]���r_�?%�?1��E�y�#�=A.mW{{�m�),�������F�0�ڍ׃�W�臘\.��{�0/T�$�?S���x��p�{hxW�M���CLO�=W���$Ͼ��e�4�gh}H<EC0�u:��6}��2qr�-��E���?q;Ƈ�vfUJW9��~��U��y��A����mftf	;p�b�c�kW�9!fP0D�`������w�0Ԥ�<B����u}[=��Bjbu�~��TY��Rw�K,���mh�����J�����Y��1�9��?���J�j%�L1����һ�6���w���A��H��ȝ�t/���-�K���0M<tMwEQ��$N�(h<cp�M��M���dQ��n��.u�,�ݼ�A�^>��mޝ{zj���20c{,�F!v]T���f|�3L^�bӊ`"I�8^��G91�PJ��S��Ԅ�.e����1�>��]�D�1�c�n���������dF��,fp��q8�wb���O2��84-���yX�k�B�[��Ի�1{"��*h���u3
��#4�2z��>��8��m�Al�,a���K%�az'w�(_8��5&GVU��~��!��[�w�}n|]��O���ż�Q��R����#���q�VM˛R#�4����w�:z�ܤG�������0�j��h ��P�;�+�Y�@zeo�{�8?��gED�2�t�1N��F>jC\�Wy�#����.h�PfC���#f\�y���q�i��vo�����j]8g��M1i�t��Y\�Xd���81J�7�O=�i����of�b�t`2M7P��gu�?5��.���y�Q��+��S�*�����˅�C{c(�m�A���IV����$�<����^��-���b:�C�Y^b40K�)��]
:�K�\��8�XSd�����J��X���7�VO��}��Vǚ�Gm�����g��$�F@��]��g4�[M�vk���#���t�?c(�7�c�9Ii�x�Uw�ypt)��#V�Z�P6u��u�ف�E`P|�~�F$�A���Yf)фjU"W�� �����]l�Ol�j����)mG�q���A� P�	��<�g׺%�z>�E�.� xH�m�?����'70+DVl�D�d\�%h7�{)���H��h'w��^[��w���e&$���2d�����L�pt��s�͂���$'IYN�ɹ^���nD���h��r`tr�B�책f<�`�b'���L��~>�ݿ�ˀ���'�s��Ү�"��k3s�RsN\f�)�nJ+ɦa��4Џ�迢E�W?��ɕ�����_��S*^�F\c#��+��rq$>W���G�|vǉ��R�JR�s��QOcXؿ/0t����oD���'�^W�&2Ҿ՛l��_��X!ȕ���:��DUJ�5Gs6�g�m�þU`/ɓ�b;�^@�J�w�Kw�7�?=��.�ю5M���ᔧ��T�F"L�q��X��] ����O��R�L�w (�&Ĩe�8Sh)#a�)��>��k|�4���t�u`4ڻ]���	O���:n03k�f+�ˁ�
ט� ^�d��Aan�Nq�\���3�$eaG]��{�Ge7���$�Jg��~<z�]�Ɨ���Q5?�M��z��+����!�=�O��l�cu��9���r��n7�������I��QBy�?�����e�����=L����?|Q�Mz�X����*�=-�A,�T�V;$���A�+�f@j&3ϖ`H����5i[����_��S��k�Tj��iw>la�U5��$"B�	c�BRV�v��as��qp��˳�v8e����I�������^��ڽ�h��= �}S��7�O�Y�rkB�T�󩉁M�7���Q�k�F�-q�9�K��҇zX�, c�g�
Ԁ�p��}Ǯt%c�e�����u
�r�Yz�&X�������yQ~{��Ŕ�b�Aס�@Ӭ[ա9:ů��i�8�Ȯ�(��Y��$mt�(������A l[�?�<�Tp���
|�^ް:y�$�hܝ��"z�O�EeJ���J���b^���R���Ȭq�Nu����B_��
�9���(O�A�
�c�*\�b.�Ǉ����G���].SWl慩J��
U@�*\S~��B ��z5�3*<���\�;h�J=�3`rV�ܣ7��(��O�#q���b�s���(��XN��жh La�
j�O3�j��j�K��v�Z��vX�	=�qٜt��#�`�����J��a��/�T�`��E�G�ٮ,�F5�e��W/�*1dͬ�?\~#� ik�@t$,��*�o���YmGƔ�y��B�S�X����7Q�!��p�BT�4Vq�I*f.#-�/��j�7B]�����"����7n��P���L�� �8\y3�y9��^�6p�%k�I&�[#oD�N���m������RU1M�n�d�_E0�Q�}�Ѩ�E��9@��;�^~���|����9M���Wy������G���g8#� �41�t�B��!�����c7�����~e6�R�{*f�`�/�n�؝��C��������)�<�Y�.����9�6�^��g0�iVR>����)f�9(�|��~�r�I��f$?y�?{�H�D���W���h��ǂA$�q��i�Ҧ�:X�ʢ�0������ �pV~��xJn��Ot=�S��Ow�f��g�ϗ�/_���r���������.���Cpu7�q'}�_NT�$�tm{����T� G���U�[���)�iq�|p�%p�R�Nq77�?l���v�[CP,��Re2!n���U?��G@�8K���=Fq/jGFW���+�����#���-�����9H+��5�D�3���#ީ�cs:���\Y���G�����:����pp�Pû���mȚk��}R�]q�Rr9�0�k�2/��ĴWBE,>v^��	�F��&A���pZ�g�I'9���9WD!�ԑ?����)߈O��Rf$_�H�vz,˃�t��`�W�K�d���9�W��ĶS02w�D��1?AW�?n�5�TŻ>Zp]���Ŝ��6F�j��<�l)�6��Rn�!��c~G�V�&��j�M���6i��<4��#�o��=�Ӵz!\)��ÍrlYq��{�rU��C� ����s�����`�0\�$��/�p��K�R�/^�܈l��Or�^X?���oFm���eh�������X� j�� z��M��u�U�ƙ̚'�"K�v��Q��͟�[�$�MX��ݍ:8o�^�1�
����`�>m�%��i����*Q�K�Vh0��Q��Zڻi���W���R;��r|�={����t�Kb�?*(LWEp����H�_E�z�}ˏ6��8�a�0a[%�7�e�]?;�|�$�����I+�D��M7G�z��nS�ҥ�?,��3�x�����KQ�;��?��w<��Z�W^��0N%G��'��HOvX�f�Z��DM+��xAv(�j`�4���7������1^Sy/��.�u*HMU��ۖ�1a�lګΙ��HӲ���IG��*����� ��M?k�'�(p��/�~Yޫ7q`M��c�qe]A��q, 8�C̷#5Br��֮�s�Q���׈+��"��m-�E�P�e��+!���}�\��肦 �(���L�� [=h}b����辻T0�Vh��N�mtI�q�s��k�R\�\��v�P��+���/(Kt��ڷ��T��}�FE����j��Q�
���.�����`�G�z�>�\�N�p�[��]��}½}����J�ͅq����l{�Va_��W[K޲^%��V<��Ϥ�%�8��,-"��73
�M�ؙ��|a����d��C�`�-��)c����ӥL:ܝo�"���`p�7N�SaJ�O�ЊP�`��$���м������T����C��иO՞�!h�pOÆ K��w���9e��M�~<o��.�C�=�\s}�_e���9�H�F#]|���:��hl��Y�ܸ���mpR|�H�-��B6�)�L��gs&B�G/z����\��-��(�SU�?�n��k�.��!X�A_�+��ء�{���ug;7^��U#�!�V����U[ �9��`G`i{�{R����U:Y�S�3��Ԡ���u����v��%�xk$����Y�����ˑ"3���.u§����R�_�uq��C���_O��շa�� u�X��&쒦J�U�PW@������0��Ǧn���nV��3ž#�tq� q@(/|�`^e�,��H ��Q2���0�xAg��{>�޽
�T��`�%<i	Q��ȭ~ �s�)ɭU���{~��e����l�C~.mg\���N�5��b)f�B'�W����]/ߎD�Я�R&|�B��ԁ�{�`�t��2��O���G<�Jf��0��`T��%����_�3j�3�8K2����g��>��[�e�p_h����C��~��O��3�d�c&I�*|���7��D�e�`E�V!f����i�Ie���U�� %�D�&��!���b��(|�����_��M��^M�GIze��٬��۶��/��S}c|�]�����C�a.f�	�#23~Ti�<�R9�+nY��h��eC듇!'�*�����4��x	]˚��`e�=�@<�1����G�xr���6'B���i<��1��w}Tn\'ڽ�%�{`�q�n�6�b���ݕ�Ty��*ox�U�Na �g�{�w&%d�
��BRX6�~A-�t�l6����?�t�05A+:�A�Z ?荇/,{~�	#2O���vhG��d�(�2���xZ>�'A����A�3)��z�r||�!��ީ�&��s�����W�-EH*ܷ�'Dp��G�oy�Ԫi�a�S:�`��%l"�L�uz�Z=AO0}�dLy�mF��]�rÐD�Mz����V�&1�8��t�E�?P�ĸ-M�X�E�nR}@�kUI��/�"t�=�7Z' !Ӗ�%le� {,2&�{�H+v�N��<{L�]���o��9��|���!�Vϕ���r��d�R���ټ�?�_ A���@�%�E>`�U��W���xݔtm�]�}5V����Du��p�fB7�U[#Q3vT[�װ�.�ǩ��3���xP7;oݢ:Q)o��?��C����X��>�j���A���n�_�mD�N�rH�!�8�B��2�Y@viW^ �P�������Ghq[�Ԛ�kG����W'5jə��ƥئ�]ӎ�����<�6d[���ɗ1�%�XF}a��f�|>���.ƛ��5U��"���lL�qa�+�?II��_���oQ��MI������eb�y4v>�[�4_��Y5#�@�&�:����A���?[��Xb�c�c�<ͼ��eUA��:x��@�4
�B�=�)�*-6X��X���ԕ�+�v[��3�>z=A�ª7u'��Ti�����y;�-D� �-��bQm�*bu-�8���(j_��r7�ѐ+RP<H#�5��ح��{�.|����~ӿ��?I����%��e��[3-Ryď�W�V��=��;�.-��.Ȣ{hF1�����u���Cf��Q�Ӝ�Ei��
�(��T�=/�F�}^3N3]���T|�?l�I�[�=�ϊ����>�#]��[�")	��T�ПU�l��C�h��(�������y�V�8�Ȁ�<��
+|�}�����nFO^��`��B�q��+
��������W5 ���iX�����kI�~M����g��z�;6�u5F+8C�;����U�ӧ���on���<���OŮ$��)�@W�RkQxdlQຬvR�c��"Ήx��K�kR>d��x2����)μ��m#ڜp���x��bx���yX�=����|�u��KX�_�h�^*��" �>D;E����j
�����q#�6�_��S�?�|��[^�y�F�ԕ=�3/��36�LZ��"rдN�bW�����D7��/�C�a^�[cC�Ξ�:.�1�����_\� [ mV<D�
%���rwY��;�?���X�ٶ�2y��Q9�.L��T�n}���틲w;�BM���z�*s�х%��6�cTK��H�ǝا�C<��J��X\��ԸpT"�T��sr(�"���2ZMˌ�Sp�D<�$�#��h�p���~��(��"���p"�
Du��Z��OE��`~���3�3����]a{ugL��1�ʏ�� �T�f�gb�IB�<u[����MU�K�������ڌ��R������)�jAF.j�'�*ۿcP��Q������`�I�'̭_�+�V��N|;��?%�d��>���;��qԲ �E�*U;��*�k��V�,6�;p��K�u� ��V�Cٲ�A��~QsS&nO=�d=}� �/v|-v/0X���&X�1�	�c���}�nJ[8N��z|�Woe���(,�iڟ�H|�Pq\�t��2�hF�7��=���;lg��0L��*ZDMQ.C0�m`�	4�_���nb��{T�����m�̄��±:S@���{���P(+�ϬVO2�m�*ş�u�3�%M2�q��k&H�9`U�~pg��gn"N,�8aHp�����v��(*� ��-��ޒB�ά��P �=hy���q�jK�yOqbׅ��Xys$�,�mp@�g���z/|���=��] HtJ��S1����*ׂ�D�2�DV8�__�ؘrMǄ�w�g���u����	��9�|Dł�F���~�>'ѱ�1G���{j�_���[�BX�y縗�n�-��݄�0�;��_j |jnv_mV�+t�S�fcE� #� .*��B����/<ˋt����lx[i� s��OA1K$M+9��'`r��oW��%�u�b��?�I�r;~>>H�&��5.�v�4/�]|�w\$C?,ay!���-2�D��bf[�V�gs�s����o��ϬC�%�ftF�m��}�����~��� ï��ԝ������s���N]�J�#r�&��/��م�^�^m���(_�?ڐ���-<M;(�z75���#n��u�OU䗳dv��.Ő������6��-O����ⲭ�bk[��@�F��]5�0�X��,�zH�	�2�޵���t� �1Z*�t�d=��_������J����V!�sE�r���*P��P�Z2���Vxf���8�jc�'g+R��C��,��$7C����<�4�-,,���hj���#1�S��ߨσ$�l�r��d�i��q�t��Bk�E٣��/�c�)����wK�K�}��B���]U!�Q�o����0j6�8�K�qP�7u��-醜^y*o<�ƽDww9��*g��FQ��޿߰1G�"\��u��|l]�߻1�J�x�T	(�w/\�dz5��e��=���U�w���on��t�F���{I~�tĞO9����f}<��������bȤ�o�ND��,,����2��[Oj�Џ������>�qd ˏ�5���\r��|u�&���k�vi�}�q���0��'�� ����X�S�+34�X882�#����N�I͢�������:�฾�i������U�/������ �)�6
y�P�8�jl*){<痌�J�V��G�gEKs�˝T�G�����@�7�Y U���R����4B2�ݛL�_�I'�⾯��R׎Q�,�&8�s3��H�9m����)�7�gنN��SH�-��O	�wA/a�O.�L	!�|���w7|�kzU��o#\4Vs�����|�����v�����O������PN��v��n+��^"�F����Zj`������L"A<Y�(i��{Ń��s_�\͚�΍�go���H5�!�4���JT��y�h�am��s�/�T����oG���7�"��"*@�WTf�]/�C���{�}�*���]���>��pƪtR��>	�G *p�@��qv���ʎ;m����n�%�ݙ�E��i��Bȹ�#k�tЁ-�e��#��'o-�w����ذ�A��������~� �e�`�yg���{�I�-��><�&�jLtge���/��F�-�*�����'�c��a�7{� ȑeF�n� �����i�/z����T)@����)-�G�y�#W6����j������3��y�y�G�o�Ԩ�
E#v�8>�2Q�k���[����i�Y����dQ퇄T���u ���>�\�Q���i��4�]�+��>�����y ���dLR.��*k�-0����� ?W��,�&�I��x�j�H�@BۀqnWa��*�r��мTz��.�M$^#�@>qW�`R"���1�������P��S���w!�@��gM�k���I�^�,Q�'���K�8�Nб���IO����e+<V���U��a�ސ\�~�^$Kt4Y�	���l���M��3&��`Ͽ��b��?ƴ��U���?&�^D��L��,@зK1����.S��L�kC�����v��� �ڶ���bK�l�m�ÿ*]=�����^t��Ck7�N>{�Q��p�l��E��8O^@w���`ò�-�v��i�|��n�J0N�[��>�(V9B�<M"}�6&-�ݙ' "=��i���4��^GdWDB������:5{z��������2Z�Q-�׭n�A�Q�:ǹ�(�~�{�n⭩m�gS"%�Zya.��r�)/E���+}R�)�����gM���'��s�ј���$���/�8��(�
�_����BZ���e�7���t>�e�e���+���h�r�z݌��`�F�h�wD[�f��$�����o�F�[H��G
4���fQL��sͮ�~�����/-E�f��{<���ں�li[���=�J���ضM�D(�����Bv�t��t>Bob�׬���y�����4qp ��ǉ��Á#���΢5k��vxH�lT�R��d!R�B3����n~ �K-{�Y �� �̜��[A��]{B�:�KT�(XE�:X�QfT���:���]�(m�RH����SsG����Z�e�F��y�2�H�G��	x�YF.��:IZ�Le��I�N�P����d��c����9��<�ңx=�� �~��\��ᘈ��D��@���]��{<b�	�󭻡#G��ʎ���A������+���b��Zs�ԦOdby�*zK��&��!�#'1
��䟹��:`^yģvں+�m�� &�3�	]4�5q�N���lJ"$�,����' N���_1�wý��2�Z2�ٱt�v �tK�IE�4u�1�Nzc�oH�\����D`�I<�"�����8���l�L�wU&vm�XV�{3�`a����!��U�WݰWv>��N=^'x����O�[�����I���KX�w��̙��s�T)w�+�$劊z�dE��%&3�\+���<�8��u�-�x��Oَ�㩖���
�nl��τ�M[ʉ9� <�9��?�ӫ3Q�҄cx�00��r��,�>Z�h!go ��Da�=�xv��K*��V
_�����(M₂�q�IN9�*�9s�')A�&÷kmte=�*��l	`�5 /N�+7��KB����h��#7+)���2�ܙ�!��TgwȄ{�m�O�O�~�H��0�����u܅���::���'��X�D����E�%��"�H�@j��L�:��Џ�*�V�n��n��9��p?��gl��LV�WN�yE�!���t7�>/�u��r�q#��\��\�뱡��e>���j�J[�^6�W#��x���5\��1���b��b;N�k�H<�Qd�&U@D�7�#��;3�m�yX��߂A;��9܄pl�����+��]��k�]��_��&t&<���O[��'V0rt2�oz�~�ܖ�.�9c��WQ�f�+<��}����������K����]���2�q�^P�YK�;��x܎�������f\˭�����(a�a�r)�O��C_ά6Ӎ��(9��J��ov�G!��ܵ~�,(���C0\�U�~Q^Gܑ��]*��X|_�\����x��O�+�;����=F�x���Lr �����j���p��,���۝y�h�
q��1�� �XN#7?:K�M��T��s8���
�3
J��FT��6GnAR׶Va��봥p��$��
y���XUt���8�_V����ϝJ��+Qj'��?4�%H�У���Zi��|)*B_C����P�`kZdC�B?C��(���x`��k�P��X�9� g/4�^�!��?Z�eP=�®����@\����pF�������a='�b<�P�r�W�r�\�� �%OU%�h���
�p�x2aى��?���LhW�		)G� _��R0�[�Ss�� `N�rV3��GE��/��\!�솦u �$"����/�v�D�r��^>|T�O�z܊#� �	@�@�pa�pEp������Emm|�@nq�G�*�T@��)K�aq���F��*����(�(#��y�QJ�}�o�xc��3xTZ֊�5�fQ�Gt)����
HwuՆ��^�'���,��U`����e��[,�}V��iK�;�8ьo���#��&���F��na+S�z'���1�Y܃C�d�2�[~�C����O����g.Y{�ӆ"U号�-%XT�{��<2�n'��E�9�o�g�
����!ުH��q�!=�r�V%��%�B���ڌ��͚���5��ƛn:�⸫�q��¡��(鳡�m0󹝣�G��/hQj��1[�A`2�Т\Q� tr��!$�#��yQ�AH@E,%LR�!����0:w܌�X���O�l�p,�0����^3	��'�?�x���_�8�mu�?�m���o���'�N<��__�Á2�NZ��ɾ[I���,6=���0S�p^�XB
�pm�Uz�`M��x8x��7Ea[�@���Y��+�R%��������b�v0�q������p͑l���
!.��㗾sDE�N.qy���4��nY=>�1kl{�=����|#�<8x���iY�?�U)w3��g%M�Y��o t���t�(z�F����5��AhmÌ?�ڴ5t�v�j�HY��A`$1�ثom �p#�	��dK��,����A[vJ�(��b�ϻ����b���u�j,P��C��([��k��3�H�@S,��ڻ��+�)B�mL i����=���nr�9U��[ǆ�y<���X]��=� j%��4��0�䈴�T�i!$��B׀JK\��i��l7+�K[�358(f�}��L?�یW�C��ιʃ�m4Ni�_�;_E�9���g!a�O�I��
#u�s�*�:���c�lML��e�Ѯf��Y�E
 ����Z�!	�=R	�y�	����'�&���%p��+v@�ȅh`�Γ��Y \EGC�Z;�4Y
xK�-4>司��?8/˃^��]�N�K�I���Fm����}'F��2|�D��q�,Mq�m����C���)�`c�ӾSB�E[Z%Zj�i����Sا�� ���EF�Ylw�Er��0�4���`�3m��:*ц��L������u�]ծ�.���xIh�f��g�+ح���n���ڜYY؈4a�ɚwË����=��BQG�Os��-tvv@�Ӏ�M{a>6K��u9�Kg2|6r���"I�G��������f�'���������Ĭ���Ͽ�L+J����)Q$#C5�y[�,fac��ģ��y�(�4��e�O�Z�8���XBe�B>��4$_�U�(�J��տ�G&~��#*t��}�^;�J��}D�r^�x�O�g��A:4=�֤�I�P��ɡ�@>"Q���	��D ��լ��� �
,�ʶ�_��>�'�����Po�z૤�:��O)��y<$R�^$Fs�ǁ�����@0m�v���<	�9Qy�����+}3���Q����Us1�3�����0Ø*6��i$E���z�\T:;N�ѽ���Ǜ�j�d���k�l��Kb{���L�E
]����k=,�m%�dW�D��7}f��k������j���̩P���$�=_.�G���A�a�A���B���E>x�5��F���b���ǐ���N����<�������|ԑ#9����ּ�6G%�S1)Q~W�O�`�;�pU�Xǟ�˱���׌��W�5;��ʂ�]z! �Ƶ�~n� sأ�� ��)7� �F:*)�� ��k/o0�%Խ��	4�
)z�v)v�����b��.My��g��tm�LZݐ�s������Be<iذ`a�� M.e���|X�x������S�>�$�����P˳3dӰi���ǟ9��0y���R6\ϔcfz���Ho:�c��}��F��38%�arƆ6@"`�n86yP������-������ �o��7�\��f�՘��2�c؝����yL�¦��ě���1�~ ��QA��Q��
���q}��"���2'p��I�1K��?�\�ǁ��>����s�Ƌ��ݓ�r�e>���h��Z�u�� i�wTc�re~���/������$D52�n����]|�Wz\�U��F��\���l��v���\����0�������1o���Ls%\�Z�ә�vN6��Y`�-�TUZ}���7)��x�.�;ѵ��+�d���4b4��NH���J�^�%]��|@m\Q���4�Ҏs�YJ�&�y h�r�$?����^��.'&܌�F�P���A���,�p3�,�s�&�㦱}��0] kn���H��t��Am�۱g�F�<(ʱL2�� �;�Z�#����Å��ʸe�|r�#nQ�|sh��(�OM�@o���y�E��0,Gr��s �v�#��f��
��C�p<
I��i^QE;�U��g�1z^P�]Mjt�{���x��c������>���%;�C����JH�hx*S ��������K� �?�"C;I�rD�f�B�4��Z?�aMw=�GY,��=3�]�Y�J趀���Q���pw��$ ��8r��	�����p̮�`T�>F*#==��m*�ǝ�`��3ۑ��dY� Qd_��H�/y�'��/ X�P#w�,㤭�CZ���g*�͛��;�SQ7ƍV��>& �o~3LߗlP���s�'���,��
ͨu�i��и��'��*N淎T����-���,�<��_����(旺@�ޔt�*Y�H����7�mn�cn�ZO0P��T�0�M�&�%@�V�Si+��c����!�T���ҳb��>�7�*�Qy���۸��;��Q�E8�+�{��r=���&�1뇍����5]�ޒ����{\�P8�U�'h�V��O�Y�i�~���ůܼ?u������D	�|Eo�����;�B���'��lx IXu��<?�O���~`��/��T�;H����u�$�N7�O����i��!��4��
gՖ��ǟ��Q��Ȫ��:	u���x��*� ���r��6�5�!3`yk�Vw��5��n	d�ms�Hs.D�����U��f�_�T���~�NU.J4���q���w<�/d�F�'��?��s��W���X��{��k�f���U�C8'�()���0Ϙ���Q_�����K��P�}ƻ
�8~��5��X3W7,��+�wF��{�[�5��G��� ��|��8u��ڀ�:A6�&dWPlr��|>�1Q���s�:hu�.�OSfh6�>��t�M:�KH2/��Jg*�W���?��0n��T��oE�.���&����c�@�RQ}���l8�L�WS�� �G���[ ���J���n�P?ԠG�PrUf��B ��V���x�`�،d�IU����4{I (^;���h�f���0%���$��`�z(��J>�;�$�-NB�^�xHJ�����GW
c�q���|�PE�`n���ތ���H�������� =��*���#�������O�F'�A�4�xܾ��$���dO�]3 ��	jy!R�}��eQ�/�L1���Hs}X%���-�PВȢ5���It�R�GQ����V���c�z����)5�PAtliv�q翪C�k���<��"����Za��/�q�!b'!>�̪���CQ?r�=�߮�A?�q���\��^bg��a�>Xl��UV�A�;Ɖ��ѱ�D�R�+=X��b��7�-��P�X��� ��-+3m����T
�����g���O��ˎV�N�F*f��FA�s �
�J�ݛ�aq�I��:��}�%t��|����	H=�g(�S6T�-�l���!�$�As��?x��3W�qv�jM�M��O�I�p�L�/��(�+�0��.-��8�(N+��[\��u#�ḓ5XpN���C^��0n����KCn3����(S�?C9oQv��h��]�e� ǋ��y�u���:Ul�qYMI35|��}�@�TC�s��u�fLy����Qк��N3�iև|���O�C؃��w#B��}�݋1y�Uգ��[x�S)<�C���E���/���!�5�t�H����¼�����/��}Ց d*|v��d`[ |{���э &�G�W���	.����A�Zt�|�T`�D�Rr>��>���'s�zy뵠@���P3K�b}�
Mk]zE>@�M���> �$(@��$-���%��n��[�d5�1���./�$_���3'
����`�k�V/�[��vC9����Q!��u��#�IG&6��'"S$�!�5��t�ȡ��Wy^f�S�$ͧK�f���g�������֔�\ki��i�^E���T�20R���nG��l�JQ;��Ѕ��I��	���gk3R������j������Z���;�d�έ�KG*�b�i,����fU0�n/�����wu}��C'��Q���� ��;/^�OL`��4r?�=ϩRe����4�%� z�,>������ɿJ�=_V ���\����:\~\HA���~	.%v�����<i]o]�a��7�Q]I4�i8؝1Vƍ5*���nֿ��uݜNq�&��t��
z�AX[��6f���!�9���,Q�c�v+��ZLQs�p;F�]
�zvG�s#Ш���!jϧH�v��j?h
���ho�?9�"��#�sE�8��\]�E}sx��	V� L�߆'Km)���.���-eRɬJ#e�@�|�ם�KGr+p!Bm�6����*�0w��
�X1�F+���fQ���޽���sPeD.̆��+�x�:�q�&�ZyK��et��(����N7��6�*��A}�;c(o�a[tߡ�BW�Cr�����y��@�1�o��G��Sl����ͅu:��ȼV�}u������L��yT�������pt�c�t���7�{+���'��#����Y��.x�@��h�~Ѿx40���ěE�����$>�8�>A\FkG���4����ӈf�-��-�fE�`�8Sɉh��X}5�(y���Q�L��`)I_p���.@X6�<�(ҁ��W����"m�!tMn㏪3�V�>�����-q��H<c�F;jq��E�1#��n�@q�^��՘Z�fEմ�C�h||��O��
��q�;F���c��&<F�
�.�p7(�CVo�$4�u���*�+� C�xLѓ1��A�P�*��tLS=%$E}Pާw\g,&�|��T��K3�!�J�ez����2��wf��%�=漼�y;+3�9�tA��Жk���E3 ���6�0�qX�C ��{W�p��I:�+g�I�w�n4�uNw�3C���X~ŋ �/sT��P���|v>&�l��R�}�S2�� �LZ������1�x:��bF�:��B�}��8{��K����]�BG��
v����6�Ry��#��\,�ѩ��]Ӛ���"E���8겧�<~2������MRϔvQ�#�VzJ�L5���(˾�XG*���Uё3��Y�B�Cvi t�zӛ�)�k%�̰d�o���fϴJ"���vV��tX�KMk�9�f���(�=��'S�a]BD�2"����;!`��;p����&	J����ڟ}���Gq��c'��e�gYyk�8���˂�^������yrP���_��q� ��bv�8 ە(㟌��	r��?��L��|.�2Q�<𯂅k������6i��hȮ�,xu�AM���t�Q�<��fM)Q�2y��S��Q �jd�����G�0��̙�yF)���𩉆jn���$�8O�qwX�A�z�2����V�+<�ma�NN�
հ)�C�"�,U�#��ו��6�ND����N�{��w��J����Xsi�o�,�D�#�v�82;� �>�T��\4�	�q0�D,ʽ�}�@r�/ePN :,�ɺT�Nh��	_������s����R�ems�.mR:�&��v���h���J���?ho���f��@:��KI-�]qXu~�ZH��������S��qi3�
���"�=a�(��w;�y�g�� N~{?y�  ܭ6UBD%��@�i�|�TJ� �P)�-gy5x�~6s�y5�9�ĳ�jV����p+���>���J��X�?���{ ��N���-^!/�*�'@���ŃQ���y��cF�H	���rA�t��c(��%\��=���P�?ߪ]H�N���^Z�إ�{ �a���R���-y3&Ez���z{�B��.����$��^�-
�!#��c�f����&�Y[����~���7��ۅ>A!r⻠�M�f����>�F����5T�Mo#̵*��ޖ��'�(�k�~���4��� Պ��B��@�����cl$>i[6�H�9�"DD�[�'m" }Ѷ:;XV�{4u��b[�q��r�U���DL`�G�"��)��|J�g��0��W�_�S@ �Q\���"V��a�ba��`�M1A�=dx)��w��+��݊(��炈��fsD��o��F����x�'1{�[�1Xpw�������#=�v��x�"(j�0׭�=�0���,;S�QZaI�5�` ��AP}��RS�G���X��Y��<}B4J:C%En�D�`-X��g�тY������h*ϐ�B��hO?L��P��g$��Φ�)���z����������(��p�%�X�
=�����q����J��G�Զ��.�S_θN�wU?W �
Q��C�p���l��)	��=hľd,��%o�`�S<�
�p>��+���W0����<�쒟�Q�$@=t�,��
���}k�1�aX30�c�'�����VyEB�><�p#�h���3�N_� 5�q;w��p����_ʖ`�B�/��<�T(��R�N;*��㹰
\Q��^:{g������D�8O���R��4f�O�J9�!wO�߲ބK��\�,�ZƸ�,���Ys�׼t�?
.������X,��ԕ�u��.��Q��yq�+�;�Ob�9.��k䜙�`Gΐ�8Q��蜄~�\�K�A�;_�n]SIc|���~�yh��9��2�6�pڻ�d��)�5? �J�>�!����D�5Y.3`���ͅl�N����͡�j�# ��#B-z:ߍ͑"�7ͤ���9��,����."=���=��g��J������$x����|Ed+�3�D
�#U1�t���A��*�~C�5HQ�E0t�O���_NYL۪� ´3]�20�y�`�U����޲�0�߯;��H����ȡ_MS�H*�p�v؂�t���r-���$:�n�]�m��u�h�����r�ܽ�0w�nNq���F��`�&.�i���M-�"�K
��Y�ْ�Ο<c����F!��C)þ�;���=�^9�
Е�3�k��D��mC�ر{C���'���+0l@�	���y�y�uOl�5��o���Pȿq��VK���NU�p� 9m�!�_dD�˶]�H׈S���C���2Q*��T�C�'@�{l݆�4Z�]�/X@�_z(�Q��P!� #����i���cS�~p�Z;�y�摬����@��;j݀����~��L�\M�+LB0���;������Ψ��@-'2�U��@C+���?{ⷨ?���3��a���H,2�������y�;��o�U��Od̆�vSD#�L��&��c��ͧ
�N-�G�H<S���_6)�_�pnX�+55�J�:� �u�)
;7��-��OB��d[�����f����'��ꑫ
?>�[c�_�|��Yw�*�0CУ���=��ͻ�c�0��c��.�V�ɷ(�8�q�)�7�K7~�%�f�*��⚉�h؜��E3�E2��v����5ZW�V�[�p���DǪ�SL\�k��)����>�`Y�sJ�dtp
c������yW��1L*�z$��Д=�"PH�ak���{^�:���\�Ɉ�$Y?�3�n���P�e��A�ؾ�9is��T͛��d*H������X�ԕu��4��~�Ib�=sO<�7�^���PZh��ĄOP�܍i���t��� �A`���2ѿW�z0��Ƿ��N���ש�j<o��
���*���������{V}�K<�m�B������U�n���۲��L�)b���W�RW���#�8���{��ՄI���|�=�T�n��ۯ���]��`0�+�Z��� ���!����M�θ��gM�k�O@��t�»�	ܽ�)�A͉���"�JN9��~u��W�%���4,x����3U�(�P�%����g���w�+3t䛷��|�$�v��Y=ΙL��x[��s���*d}g�L̞����v�{C�Ǵ�J�n�����������a�9���WIi�M����nV�c��������l��]�ʕ�h��KW���ո�dcXX��viVg��M�eG���.�E����Ѝ��=�vF��Oڤ&6S[�8�~�+�����8�s�3�" �:�����,_� {P�����0ZB�4��$3[Zf!D|JaG{���D;�sc�Q��,Hw�7��TQb���A����S��H���(�H����uЭ��%qPi[�Sv�!���!������W���7,i����/�T� >l���2�{@)b�i4l��q��䗔-���ˡ���pM~�F�ҁ�|}�Ʒ���4�z�M���	6T�g���+ʱ9z]g̱�H[�S��G����W��m��R�v�xI�׆�g7�VC�@�w�~�	���}����A�H�,�,LI���ByF���g̀��!�R����v��ln埆=�T1�T~�����K�L0�M$�Lq�7ւK�x6 -��g�_"��၎<^�@�@A{[��qt�	�tN��K��E�e�N���5d���4���O����=���n�CLil:�a^d6�`��CGl��Ya������]]��z�n�:�#nK�+rj#϶?	x&ə&L��њ�=ο����jGYv�&��v�jŋ}ٵܪ'!��ې�(�)�"x�<`*bN�um7mX���#p�!Tʆ4R�2m5���ۃNbπʣ��+�ً���{�ˋJ��Gg;��`d.���H�#%����.N�U��1�i�]�i�&۱���K-z��4�yx��x��;�Ʒ�4�`O3��U�n���l[�_���׭����;	��� f�
(��kU=>xc_�E�%Ü�sz2]�U`W���)�f"�BCWe�.�b1IzV[�{�h/���,�c�u����y�C���"~����I�.����G+"�.���<=!�݀������m+<gON�k�w�"���9��$�@78�RUT�}��g�Ʀb�K�2&ݍ'"�P68��q��e��¡8"���}�]�Ǧ���Ĕ�a�-%�0�0��L�0�W�qBZ_W������;� �"<�2�'����V�=�R@�z��U��H�t|�22�<Vf}K[�%	L��P�S���(?����Q���I,�)�\�m=ťO�G��=*$��8}�
�S�e��Z��0�m'=�<K�f����f�.?D��N�|��Qbu� z�}����\�A��P�o:	F�ьāP�|`1R6}&Wg2��T`=@�j��9ī��� �l[P�+������Ue(�k�����|�T���;K��aB�r�̨	���Y$�Ǝ��i���:@���z��_:�>ڥ��K`��[��U��'%�8%��=.����+�A�d��_	�Ń?�f��X�}�*�K0���/�1̃d
��Dj��e-uT���ߏ���N�fE��T�3�<�r��;B�k�;�8���u����Ð��@�ӟfN�%ƫp���$�oG6��HՐ����ٽ��QNU�9�&I+�#=�)ޠ�>����}�oR%n����m=���q�aΞu�C�J5�8� ����6b�X����Sۺ��,X_�?(��o��1�.A��.F+�I�G>�Kh�ڞKk;O���=��.yc�	�" ����M.���+���5?�e��\#1��2�&W���_���^Ո@خ]a2����Qb�܅`E�~�+���x>�v�ڒ�֭�S�Fn�AՂ ��^*����Y,2��=�0��f�ky��џ|W�-�10��%��c6$�����送�������Әm@� ����>��o��O���q_=[Ps�9ş�R��
 ~����z���tNjS�*"��^[���}���Z�sq˶I���~��}���iOQA��X�u�� ��'����X#I�d�n	�V���|�[+>�ƹ�V
��䤣�J��h��ux\�4��{M�ȿ5�@�G<�Z+�e���]��F��D���Sݜ}M6�Y_�f��H<�2�Ze��l}i#��e4���� �͊�3����q�o���U���<�v��V=>t^� 1�9D`wn�1F�z�`wh|�u����{G�4|�5XTp���rx����d�r`~^�����?�M�0�(�F�_'�ZZM�G��ڔB�i� � ��n��Ucq�.��'%�#*&`�wZGx�䆟�\� �a��>�#��RĢ�..��r^��<�{��+�� ��K%��_$PuE�&0�B�=F�|�o: �I
O&#L�jLMa]{�(��.�n,�~�a�Ǹ���ƛr����ZjldeC� ��9hX5q���@���(�6�h�hu�ei�J�2��C��E�O�C��\\����v>$aSZ#��&�#̞���"|Q���2�b��T�$X���|�DRhL6���Ժ�}9F���<�{�1����s'+|���#�xg�B��M�Ovt�֥>u6kY���
��@��`o; �����?�^}[Z�m����=�
p��;��^>j�(f��$� e���r�-���$����I�qO����/r˘������(�E�*0֨��i�5e��TK�XEt<�D�f_��<	l�H�����t+�w�*�jN��x��IF�`Q�x��O����GjqP8@G6�Uz� v�Њa:�>�3L!R�Nt���˿�3�:���;9mU@c��n����g�y	"d��q$�i'w��@��fyU���`��ݗ4�
��DYC�$DOC�sP���c�A�y�8Y`g��ｓ�Dí�4��+Jo�EzT"֢���!�o���?r�[ۀJ��,����Nx�]�|Z?�s箙n�6h6�s~i�P)�q�O`cd�i_�X��8wtz`ĖD�Rx�ң��I�	�,6���l�.e�w�Z�X���_@AP��-K�)�\�6�l/U�}h���P���.���b!W}[7Ϫ54��zGa��2��գ���4�;[!�z� 29��3��ሕ�sF4����zM�ۈP��T��`��̖�uh��?3��(����E옉�i�*6�����
�&����ύbfA��
�(�q#�� մ��0���)YΩ@���,B�)�|���,F^_رV���h�=��r��^��̴����`�ѳ���Nk�̣`�/":�&,d0��ҙ�����"�u��%N�dǕ�R���F�v�K��p/7��&�xwY��{�&D	�o?��ڦ3l�X`Ӱ�3�n�Vu��d�����,��n�_U\Wv�eBj@I�£���
��[Q*���F�h�3�}�������v�L������܃yL*|��m�Ɛ2%y�nNғ�J��| ���PVN�ɶE;^����%���X��	��cYz�*+�ҷA��PD��A�0֩���S�a���zѨ��Q`��3el��U�_�l�"�-�ѕ���$7���~���>� ��?����6�8���7�l�����7�H���u)��r�����Q޺s����vSw�j�� i
�U]���޴I�f�E�m͍��}Z��-�aK�ʣ���^bm6�r��ܮ솨�[�yd��t����[vp���V��8S�bU�N�g���h�3lo�����U�8Z,<�-Z���N�8���5Ӟ���7��(]Bx�zu�d��;��\;X�@->,�y~kbgF
���!���[��W���,�Zi������5�8�lcbP��Ê��>��0��4���}0}ƝB2�-��iNbn�U���J|��eI�� �����rPȝ�����#5_#�̉1�h$C�j��h �N�g�j���iC��y�#�i��~��zЙ^��l��t{3����="��/�Rk�l�V�����{�P�����؈i824!|?�Y��nՏF��-�a�V�89_&C!9Ũ��=�Υ�RG��ce�ְ�ƞ�s�y���n����"����?Z9L����C]R*������P������R�3��*ؼ��@�0'����� 20�C �$f�Ys�X�eKf�xI$r聕n��4�qK�5ci�����6���)q�;DHM����Ӑ�T��gP����6�ٖ<��3��'�,���n��Y1�.���:qX���+��(����'�)��e�^f����s�a(�ҹ��׽����sG��͹B�[Ej 2�M����Ѡ��:�$�|���UE���*�9t����:���+x��C(��x�����q8���������}=r��M��E��m�{k�
P�$����CldSr�5��!����b�S�r�d	x;�z�l��Xom�Хb
���3q����6�}�7[��")%��i7J�|�.�2$��V�4q����)��*/{��� ��Q�%H���'4M��Ê�Y�Z+E)�b�֘Sm���9KSs�����
8�!5\�<&1(;Rk"fn����h(aj�����8��F{��߹R'��oE#����J�s�c��pò;��_�XlF9���>H*�ĈT�c��$fE��H�J�l�Wv��4/��E�;73hS�܅'2�7:~�̨n�]��o�����IMO}� Ԩ�0 a|�nR:ö\СB��Z��F\q�%̓���e��2�q��ܣ�Nªp���ߝ(Gq5� �K9�
O���T�3��y&��x;H�vX9�fw �>`{�2���/�6hxf}�����*�G�΋g��S!-�'���a��|(�P�;��WL�����%{��������֢�L�Ֆu�aow�����q>�E�V|Ih����Q:Åz7�i>K��	E�Ң���$7tS�B#t��ք�Z���3Q1���������z�Kh�rr�]�@�K�*:�E����W�'�C�o	�a��޾Q��y�2��P^��|��"�6��-�H�΁]���?yr��6].�A�(�x�S�\��Q�@&�jeb쮶�	`�B�\�7�}�<��^kE�3q^+L�cV�fooҬ�^�p���52s�EA�ⴻeR�j�j7���9�Q������҉�U�B�P�2=�Ldm��_t� ��:���1�7�
�*�P6sG�^�,�	TB�r"�m��J@U�Y�o
���m^|�@����Lkr�)NR����	��J;ٺE.�na����R��z�F�_��O�	t����3��V��2P��3F\�Gu1z�l�:�ziy����v��;I����AW��Q��|]m�<a��g߁�~��	w}����!"߉`�b5'tQ���?p�8��?�<*����P���b  �o��(V�#����N��4��J!�"%����T�3�:YF>������,ަ�� |W�
6�;GV�noF6�N.��i����Cl5t��C<����n�v��P%���
�n����ݻ���O������A������3@��]4qV�K0�j�^"�QA��-*>�z骝�3������%,�k�`����,�(D�E��S\kɨw�\�|��[�=�{�/��4+�ui3��c
CIe�Р���J;$0�,�G�b��@U���aЉ�0�g�0L��[��d��'�N��Ⱥ�[oS��*%?�������+���j��T�p�v���3��a�H��R]*���ˏ��D��d�ϋs���(6>��Jl���捺Da�mk���Ԙ��]�PL�_�r�[��tcb�6���2n3<"Ʀ-��
�.�ۂ����7P��8i���L�-c+��6=:�K��g�[��fQ:T�"u�v�)B��+��Sa�t��@�8�����tPs
��0�oPÀ��]�e�<�ڣuvD{�Tmo��`I��"Ӓ���p���Àl�N-�����)	�ף#��$��%�k=��v�A�'j�7i:h$���~��N�����.�"f��gj�s�E+jU�_F��;AM]K�@��MX�^"��	���8�,�,yY\����`�:~��vx��9[A*�#�҄�?��T]����L�Om�_m�A���z���@��l�.����Q��M����Db';t(��J������w��hx�i�2���]�$R�E�h�ΈD���<:'�O�ڊ[Q�Mf�����V:�P���<U�"c� ��]��W��Ƴ�-�k�Q�Nu�"�������P�Ψ�r$���Oh^�+,G_���_
�O������ӛ$�t���ݐ�"���:���ؿ�3Q���$�)H�Ti-KP�,�\�2Lb,�M#D��U�Q?��%�<`�\�˚�[�`�}��U�J"����ܟrx;���/\�����x��/���/�W2�I���i�`n�_�cWK7zqk�*h#DSQ�ڀ�
�c|RR��zN&��	/L�2B�2]�L�9���A]��1�R�|�����a�H}��L����6?����q����.FQ}���k���r����[�ْY�7��f�+�S�����Ow�3z�n�8"�x�f�i���r�J6g��%��c.S~�/g⳻���Q��|	+�Jp���w��ڕ���	��Wg#�R�������AK�>�;l4�Lk
Ԥ�s��X}n2�Oj_�l�]�����>���9�^{T��
 ��ɜpDL�������T|�g֭*.��n�M��.��#T{7�# :G�*�!����*�/�x=2�I>�1.�!�W��D�M�jk����s���lk���a��X���,c�?�)9�Ze#M͇C	�c��FWD�}qɉ����5�.X!�\�&vP����?�t�LvG���'��z���E��(qs���NZ��5�R���>WZX]�Y���4z�d���8x�b�~ݖ�S�
 b���E8�W��K7�G�*�<c���+@�Q�����O��B#v����`��`�M9/|��t�n!�;+��.Q�c�σ�ި���ɡ�_�x*F����4���&7T�\6]�l&GFQ�_́��=˳�����
-�v��_0�g���\����ABs��Wi[[����[�Z��79U���N�*8W�9;<7�|��Z�#����[���$P��k6T�[
<o��5�����(���q�O̒�����Ǘyq�ƞŦ5\� 6su��ꓚ��H�o�OPSQ.7R����x���5 ���L|�6�})���3V��,�[�׸�x Y�,�JA7'ݷ!�.Ŀ�Zs�>wx��,���
�y�	p�N��r����,-��X��ydͽ�W��3��I�����Y0¤Cf�d2}�Xj��>1�^�墔(p��{�K1�J��\���q�5u��6,ͳ�R|���CR���`6:�>�s�~ <���G:����aStH�Wz������v��\Ǎ ��m���B��2�$2ǌ��c\�Q�.qҒd�Qi�sh�m����g��mW��U��;q�+'��;k����~g���2�[���A�Y�;'��w\�?h����3�HK���۪��1��q�閟� Ea����Օ�0))�>
���s����!�y��GT�]h�~9����p��+⡮/*�Y����'�3�R�_�h����m�����q���>��x��SC�g�??�¥�y]�{��OGQ&��W��vuNrޕa�'��ߞ��d���n:�����^T-��4N��%�i���c�d3�Wd���T�ﱵ���*YuW<�3m}�QI�?&ă���5��������X����E�W�C�~f%k�[B{u�|+r��Z�n/��M����KW�
��bu`b���Nv���j�j [#U�	�G��6��<���c�ʑ��
�O̎�$��:K{����6��p$�(���~U��@�ʷ��^����%�;��zg�K07tg):&0�5?B>F�Λ���Xu�CƮ�E�=(�eqz���l�d~Թa� Z=\	�g�@���K�l��
3��ܾ�G9|�-���w�m���˥	`��Sߟm~�̹�V�h#.qH�\_ ^s����>چ�Uл7�)*e��
l�^�+uN��+f��i2��L;���]��AW��^�n���VL�9���* 5I���9e�v�j蹳V=c��6���%�P�	�Ʌ��J�����&�Ee�����"�B��#+�%������i����ۈ�����x��t[�U���Ӡ�v �:���b���٨�ׁ���,D�]���Srl�kP�+7�"�U������ae&Uikr��{�Lg��;(}����e�{M� {�c�O���|��A��Q:�G
�S>�;@�PD���?��=ڵƺ�-Ԍ�ZA8���p�װcm�]M��1+$O�	��Vum팝��<�U�6�4�<X��p�#.f'���m~'���w3RqF/�\�)ء��x�b�q/�u�N�j��.p^NY*H���|V<��X`{N����Ҿܿ(آ�vb��:�0'�m�<� k����<��� �MN7���O�v�)��Y-DT{�j���"�<��VA�խ޹��r 5����d��D�"���@�:��K��}}���g866���Ӑ�AWec�����ﰔ��_!C���H-~��Ƴ�vU� �����"]�ù.%��2��%���v9�I�	�x���x�\����J�l���;��j�8�_*���Sz0��|�:��w]�3P&P-��sp��eko�ۻW���g:4�M �n����t蒸��h��5�2����K��D5��J`���YL��#�@�bl�j9|�%��U���D4cVU�U�7��`'����G&������#�ly�:�쬺g��I����_3�'N)*��za�r���j����ݢ�	�M̢B-����y~AI�|���{q�0@~Mn)0%��p6�2wx������[x��(v^8,mQt4t[^�S�;'_�0�}[��z?4����68;`ת|L�J�"*���D��ɟ�\
���_��ot��X;\��tĔ�2C�ȫ�`��9�U�W-glC�u����@f�chMގ�@}�Q�"��BV�/�XA�-Y=7�QK�<�W�Z��g��q��jI��	")�ri;3����\�:��.������Nr��zܷ�*��u:v(���ް�[���YufW�;�W��|�C���x)�s�.7h��~�"���oϜ�E��{�df����U2� �yp��鎣%�?�r�̶��ٰ�7p��)�Ɓzo��u��U�qH�� T9���n�:��Sv�w#'"���`�H�#h�PQ��Esv� ���u�6ђ��*���%y)nZYy/v��9R�	�X� �4�����!�`5�� ����X#���t�ϴ6�ߕ|fnA��~b^�N䢢b�`��y3w3[.\R
*atQ
g,r�%��0�Fс�N��5/���Tр]�X?׈=*�*W��M:��ʦ�Hd���y�c��	N\5��KO8§�Vn(��R�u����iiX.���{!,�Ec�� 'v��?*?TW��d�Y'�y�`���}�]`0���H�(����9$豧07��=We���e��`�Ȑ�w���{�P��5��ȣ�//�S���&�3n{�Mta����*=8�]���/�XòbR+<�4ʗ���"�R���V����+A�,�j��Eif���y\�"�@���)���dg��Ʋ��P���K�n�)ǵ�p������U��І�_�㎥T//��I���>��-�l��g$��x�9��S�D�w��/ּ>�a���cdi�/ڨ#�a���F���M̉7�׭�)�6FCP&/{���ut��l��+_n�4������Pa�g���_Л0܇5̸8��\�7�O�E$��I(� ����wL�s�#�=�� %�/|n/������5ە����Ħ�i��^��VP���bC��V��J�E;,I��L4sr�Z��c�Ip���I�kEK�<�X�-�ٹ5�\����ϯ8�P~i/\�K��^i�mљ�Vb���%�n�����ǉ�L{q�c�����O� p �Щ�J\��W�����յ�T��=L�_e���R��z�IټĢ:$N���E��莓sw�\�����%�Te���=r��M*ćR�bζ��aǼُ��@�Ѿ��b>e�H�P��{���e3ũY�--EMu�a��a,��v��N��R���60���h4�4L��*J9V�T�,�;NH�|YQ��W�����
C�b��ܤ^E�*t���h������q� YR6��/]7O�3�4�y�`g��d����񐊔u�P�E;��al�A�r=�m�Gs�ދ5�{s;�7Wj�h0�^���'�>��z���1�rcc:����im�X�i�8�t
�y&��.�٦�I<�p���22l�5�ܨ2���Y@z��\��V�Lt��SL-�Q0�T2"">uΔ���ߡ�M����CE����V̗�1m��������^�I=)�n�Ջ����c	���l���7���;�b��U2���M�^5t=�[����Z��x�x�=
#DY������qfB�ϩ� �u�����?���۰)j�S�bia�N�Qۿo�;����vM3����^5-1PEӪ'Y7t������?�DV��e�#�C ���1-H�I���o�pXSZ��?���+4��<K����� (�V)���t�mZE��͆�?�x&���+I5�/Q�C����d��,dN�x�B���<A:�4m������ QOD���ٴ�Į(`��F���̍��ղԶ����d<<u��Q;���j�ll���Ϸ�����7<&��i}]g8t	��._� �F(�-C<��T�i�qL+]:��4�9{�uiS΁W���l#���O� ���%�7%�Jg��b���A��K�(�VɎ^��5�t�>����~��#��K�w��${�^$"䉈�~��3��Kk�:�Ϗ�ư�0���g<Ed���&����n�4�?�������lv�����$��@��Hyo�We0�4�R����>Q8��S����f< ��+�d�N�*l���-v�b�Q(� �X^ZH��a�y��We��H�����8���L�<y��[��Μ41�>s��NZ�KFҍ�	�w��~X�f5y�j>��M�&�~�[fE�H�9?�
�l�h+I����6�����=�S	'�N}R+*>*~0.D|Е��hn���J��S? ���V`��W���n�
���~n�i�-g�ك�t���d�:��;�3�П��=�H�I�{���\�?~���13BV*��$���@qTp%�\&��͌|����7֝�I�,yuS�qO�6�fhQ~��\́Må��7aTs͑d7���������C:�r#�z�?J��
�B� _ ����>�k�< /q�":%�S��e5�B�P�n׆(*I�C���ݨ�v.�Y�BO7����E�	.=Qu���;{�A��37�`�G��Y�H̆�S�s߯펔T�����$�����eܛ���r�UTj��RxXR��\`��tHZ��+|:��E@���=3��@?���	ҿ]��Z��K��IAzt�ꑣ�ұB�+��m��x�4Lf�x2(���;m��_h�t����p�+��N�W�l˩ټ�������{YDl��G9Vflp�X^����qm�&E�R�G刷�l�BA,���2��-��[}ih��xGe@5i��ǖT���Ӫ���Ԙ���χ�o	1��v�T� M�s��Zއ�+�p_5BtS��E|�,i5u(��]������چy:�.���i���J�W=q�xH$lis7��j�0p1RN����1Z�s�t[S|�?�yS��z)�'
��	;5W�T�������,ݧ
�U����͹�;s%3)ls�]VP�Z��}ؕ���R�	�&�?ƅ���.���E15&�<�N��T��Bת�zu���5���z�{I���Ub���R"�_'\i�����2���]�n̓%e:�u���"�N�ņ�ExN�bꛂV��ʄ�'���#�v���]�K�������K´C!3��J}�Tf��Rs�����C��{�v�c`��l}t�#T]�����f_],���u���J0�oZ�D�!�aܡ�S�aKf@���;�o��o{p��@�Z���L�ה�&�x-d�J|F��H�jܝʷ�����1��d��r�D�l�a!!�,,.k1P�N���àR��֡����`�f��wnA�ҽ�?��):��T"��Z���@����-�g^Z;��X��j�ҶW�f%�D�rN�|@U3�u��T(�O�7^�"����`:����q�9�3��P��)ӹ����R�U�W���_x�q���4[�.p`萧 G���:���_ڲ��P$9eH�ycܭ�>� �)�Ɨ{s��[�L��t�/����!M��u6ӵX-�@�����A���	|�n�,����:�L5>^��\jQ�D/5�^�g���CG?_ť�s]z�c�h�n�b���� �t`��j6�P��Wj�.J{����zϙ�[~��Wu)��&]zb��D�YTvI̅EH�C�/�!�BƟ4_��u@�ŗ"�;���Ɠ�}* IN(�������6u�{,���,��|���;�KՓ~��n�)�ȕJVb�	� �vق�H��Q�Ѣ�.�"i��y/��&P��X���a�z�bo�Ղ�mT#=ط�޿A����%���(l�{K�>l��#��f��n��3�-Bc�PD�����f@��
�e3=��y�{G�-R�z�y�A��F-�տvG�������k�b��/^ ��=C��~L|J�<���M���s��r�-�`�_�$]W7���ұG�r0�9��/�6�|�Ne^��4�&[�C�1T�Yhi���-7������
��98M���񼭣�H�����E�Ѡ/��5v�A���]�DX��3}�WC��CZ������A��:nQ��5_@B�8wG�����ӂmԇ���&x��ƛ4�7�0C��f}b�!��m���׹Hm��xRǌ���'�W�N���C&���;�@�}ynr�p_;�:��H�"�-+3K���,��a����'J�0��&ߞ�mV<�8t��6�n��ퟅ l��GhmUb�fk��FV@�
O����u'�>W����	e8�]3�1�0��՛� ��� �\\��@�4�&��EJ�8�J�s��͜!����z�E5����IQ�+�����uJ������H����р��	�ƖJ��&�:ט4��}3E#A(?k7ꝼoI<�"ۨ������o3���m9
�Ks�=�����ch�a=z���϶��5P�C� _[�	c�`��l���z�����Ȥ[���}*U�??*����5��`����;'�Yפ5�Q����Ϳ��+]��O&M2{��Vm��0�vI�;�+��"xcBq��f��˳���Ј���^A\���nXӁR�ȳr�W�Y���D���J�oS/�j_7�>��VMi��~D<#�c�/x�b!n���GT&L��:�\v��o�P5a5���?�X"���,���g��]�;�#�c=GR�{��)��ñ�V����{��V)�&|f��J�$��?i��iÏN{�`����v ��	#�f.�>:���:�)�=�J�"��|�C�ze|���:�:PH���u)�s�s�Y'�m�����W�fT�i"鮦��w����Eo�~~��h�_������B�=&IaR���w�+U?�rw��5�7�p�崨�bկ�z��\�~�C��
{Ƶa^ڴ�O�'%BA;y0����ah2�?�{�!2�?�@�!�2`�KW�u�I�j;���� c�I\-5�����2}����&�z ���l���˛��9�Io�9�Y߅�]r�,;��I7�T�II���#�:������@z��[�Ǣ���[�]h�Oۑ���P�:f���}3j���,�=������w�J;
d-��������A.ˮՁ�Ug� ��u�C����+�C�A�z��|�3��c�ƽ����7!�c�
��-�qT��I���^k�)�@be�@_2�׽�s|ӛSj������؀�u���Ӧ�+*e�������C�쭔����;����|���Q��̷��v}��/���J�+R4������8b��	����a�`Ò1�R��5�u3���K(x���"']�~�
��sH	x3�8q�/Z�.V�����4�F�� @Vtb(�{��-\��N>���"��Uٝ���z�$f�O^������
�m�mS�!�5�l���|�� �����ޕ=����PDѦa��*~��wh*K�!g�ݺ������ ��`�!0��ۯÍg�e�YM\����#9'�Ja�.�#*�����@���w/'����hqP�7�@�����Q�]@"<��<�3k��t��2�^�bf����3����f��ݶ"z���#.
Q����-�gC��}a`�y��]�edi�fUe2J$d��f���$4�	�^]�O�����\_�y)e'=�o�@��P�p*I��+�;��B�ENIy�Z,��:7�.G�	�%�#8�-oi��A°����NOP����e�1�������H(^���!?���I�հ��M��[�ۀ��,T�Xt���P�F���g�uT��bDN��:|%�f�:��Odꃂg;&-��k��b�-y�;B�˓��}�Y�&N8�NS��8�b�J���^"ɇ�����t��@��`j�cm�H�G�ώ���Xp�ћ�͡2��uL>��?�2/�id��L��\�E��4*���w�0=���j����|љ������N���B�;ؓ��1����K)|��SV���0i�tI�r+i��
��>��gB��<��'6�V�.���a��'ɴ`pm��r]S�~z;°��[S�=~@�A��$��n�I�q�|�/O�^���Q�t|ɮe����>"e��
]ʽ�+�yZo+�B�D�z���_�F���<i��Et�TtҜb<e����&�gJ��_i�M���;�{�r��9��ӏD�=	-I=���Y9Ǔ��i��-U�ՅMK�F�N�2/���(���&M��ZE�d�ր��[��`����X�_�K;g�mG�[h{M�נ��xR�c�>�Q�z�5����1>��\*���7�{����zP��U�'	Y�J�G���+Q�Z���$;�]���B;���7ґQq��q}ȁ+ؙҁ�����[���u�f*����}M���c�w��xf��Ȋ��V�U��$��CW�)Cp�Z�M\��]=�Z��?L�
Sf���.���[PC�D��o�/vY|N?1�F���3�9F��*b�!=&�p�Bs�B�>��.G}��,��c=r�+d����66�r5^>Y�[S8)]������A�*�����Z��>2�C��+r��Yy`eA58�0C�@{���c��t�h#���P[� ��'��#Cm�~ucQj�퉔��ɖ"Ո�D1V��������H��n?J�h�|�¬S�f��!���#��{TW�i�l��p��H�`8�Q:PMs�`�!9A�F==��uI�#-�B����b�ux{!'�->�Ǎڹ�Մ�me,������t����h�oV��"ry�>��f�V�S;�����u$�� A��zpMJ�JP��>��8T)j�X�I�	�?�Ӎe�}G�
9l+�������]Kg��ÒR�3N��j�^Ϣ�t2P� KG�0���:�����w�h�"���J���E]�E��hDӂ�_t$A�T�C�'."=�i��^igI.z���p�!�orT˴S<�Yt_qb"e��c���b>��"���F��#���g���k)'{4���j5��R:,mЋܲ�����cTP�6:��I�� #�6��k��X�4q0�լ�����	Q�}��9Oo�
A$�����3�a��b.?�%;��SH�@�[�X:,`�����znj0�bH1��Z��)M����\�*\p�i���.�">E�s��>B���$	�� Y�mЂ��㓳���ã>��2�#���t^*T�|%�O�)j���k\�ٸ*d�?/ۍ*E+q�R�V�}j��?@W#�4~�w�w'6@nF�7&p'���'�j]�Ѣ��f� F����Z�I�,I�kR4鿒d^*?w�^? ����U�#�m����X�"<$���-ɚ�x<��o	��Z�-����Z� ��`�:: ��nY-����Y�M��$����y��=���;�?�<��D�}�+�q���2�.�m�s(�h�']-0%�8�����J
�rR��0���ʊ�q}�H�(���r�U+_�Qw�B�r��OpەTM��u�a��m�i�W;�of܃:��\ �x$�z�B��������h>�߽ǫ��R&H>��7P�c0�4�Ap�G�6�izB,H�=Ʉd���@�$�''�6��$��g�US}����ť��i�0�d=,�z�e�w��855߽z���7�t��.��u�����͸��,p�H4=�n�{PysaX}Y}*R;�.W�������|>���*�1��
���s*��!$��I^������7��<��`�k9�l��^EF<����j��L����.����߬�嗘��^��Ӭ��CIۘ����}h�1�)�W�&���5U9?os� ����-�hy��γ�9�W��Z�͵��ɤ�S�= N:�Z]sG��aEao���"�{��Ab�4�h��hnH%v$�gp�6C��:W�P�a��:嵊��rlmI����<�Ǣ�>m��L[)�v���'CƟ���T�e����N�0��/��t=��5��%��-{�a�x(�p��c��eOjz���r{n?�s�`�2Y2��7=�HG<2u̹ҺXƙA�K�������_����Gh������B8爆JP�_*�1}�?x}9퉺�>E�(e,pF+��b!]ha�U����B�)gG��Rx��������T� oɎ
$6�_��bP�lA�����)dI�6[�<`f��@�LXfv <N��d��<eYݹ��W"Y�7�[�=0wԗ�e~5��]^)0f/7F�N瞏���]����#%̧D)-�����ɝ��p�g��{�����8y�E��3�yqbm8ݱ���dZ�k~��j�0�m�-�,ӆ�E��Q$�ʓ���@���i�D���Tu��R��m�u��Խ*�j��
	������dS�F�4�X�)��Qn4LZY�p@�Y�1��]ؚ���xi-n±�<g�C���Y��c���(�����#Ħ8L �� �aEm��#!u?�����@���]�@����﫛|�ˑ�d=	�BBӟڹTf�aGx��>>���:�뤂?X�7P�&����l<C<(mrYw�"� ��U��X��,�.J=��O-Z�i�3` g��x�i�zPJ�z�A���B@~����s����Qt�|dqIV�H8_C�z����.�D�b���5Ah'O~�)x6_U]*6�k�޸>�|O��*��ˤ�=�-ϑ�kx��W�v7턍� ���DfEmn$�x��ȶ��a�E��I����0�
6b�Y���W]�}�i�RF�Q_�P�T��3��GY�bx޽C,}Ew �fu^EOS���g����$���X;-:�0� �%��q�B�����~Ĉ�SE�K�/!�;�ZLv�ǅ�KC�"�l^Yi�eC]'��9�l�,���[=y��"��M2Å	=�K+$��!��Ѿ �	�/	� V��
��ޭ'<�b`~D6�S&x��f|����B��ԬՈ�~,3
��"<�В�lxng~��f���z?�=�u�-F�3z}8�!�:�.��",m���FY�yA�h��/6կ���h�Rm��4+���W��ƚ���Bk�|@�tU�h�������.Tb�����9��*�
����IM�vl��a�Ռs�wp.�2�R;�=$/��|K\�x^�Q���	_qS9���p�鰆 ��E�������qbW* ؛p6���:�����?r09�.Ăyz�d1c�:��W��Ie��A��oG҂���Q�[�w�����T�Ӑ*]�"�_^?�z�p���칾��C�?�mz8���JIMM�aV�گ�+J�?����`$���Ȣ�[�kp�Eb�c�WJ ͈1��'(�B����³GV/(sŮ�:`#(%;0؜V��Ӳ�Niq�QC�a�E>�+A�>�j���0n&�w Gǔ�\��l�IŶ>><�����d�9��Xl�5#���?�:���h��K���2�;[�����l<�]����7Բ&��y�<����
�>�?1���y/l�<I�~`5	3�{}�n"�V���s?3���e����w7���a��dac�i�]��fF�����Ǔ��UlU��S�Wʱ����p���P|�ּ"����r䡱��X��p�"U�*[�J`�U�33���8�d�M }���I��O��p�h[kd�y��ϓ���080��-5�I[�`�鞇 �ēD���R�Eq4x@�g����A�4vu�t˝�`8��-�dbU�Hsd���"gaz�#�[�	�kꦑ�@qkV&Z�%%dZ�B:»�Z��)��"|J�k���F-�'y�]�#	l(ԣ�JR��L3�c�H`��4ƨ1Z�|;��X1]O�=y�^�FG8lVf/v�eզёb��zw� �䮢��F͝@�����I����"�S}��K�P�g2��܅�x�y�еs�`y�u�e��m�[0P0p�W��D�7K�\�Ѯ�,��O�.�0M�0���wc��tp�c췵����郎�>��ё�${����<��&�P{�*�|�2o�=��B��̓xc�rj�>`�{Ç�l-��En�:�8����N�ܙ�>�9��m�-;;�LR�p<�ɘnpj��K���-tDO���[d�8��zY��u�P<�xD�_f�k�a�^����\&/NU��!�/�eԾ\��K�3F�V;���.!d2��c��q%�2�t6ҝ�L~ѣ/
Nd�8�"���|�i�s{�v�E��F����[�w�4��w���B���p���y��Yy���Y�0�)4�:nִ��v��R����Zs��pW ����\�޸-z1��x�+�p�o��n���>)A��O�i]�"	��u�&�t2��%m�.==[�e\ȁ��֮�]�hF�gO)�QX�⅑}h-���qU���4�e>E��d��ˎmeR�b��%��vWMv�
�a�¨hT�-W
��"�8��Vo+x��'�}�&	ǳ�H�|�4�[B�=�۱6�忆�NΊ�v���n�'���xd���"��;~����T��4QS�꽜աi"Z7cK��*���P#-����U�ƩI�n��ν�Ϩ�KH�}��k�cp�H��!�}�ڞ�eB��Mt�w�e
~���r;U�G �I��	���v$|�wOL�#5鈐��x�k��6Xg��oe�p�r>K���EH�D�plL�$1
���x-���,�
 �q��Aq-�fX��r��
wl#w��s�뵇@b�v1 �"j��_��>���^K X�S4|{s��`����C0�/Z�7P�?Ή��λ�� ����F��LI��N��ݣ}�&>rl}?k����o�tX�n����29���̲`�	'<�7�z�jY�y�gkr��j[!�d�#�A�H/!�B�XC�O�I/���ќ{��8���э������#r2 o`��$ ��HS�����U9/&�L��z��*�G;�e�"�`Z���|LҖ�;0����������KLm�C��H"Fsf|^�E䭅E�!Y0P/�K�8�R(Ń�kUdnm'��S��d8t�I�#�BD�ZS�3]�+��6�Dy�#`����(<��y��O��5�DU���w5��:Z�� �~lJc�Qʤ�`����̨7W �sU��A�2����= ��;�r?����Ҙb_��K�>�K�ҽ�,;o�Т��c��؋#Vh��7��^����~z<:������8^E�9�N"������[V� ���y]��U'	�?t�M��8�SF��:Icj2��@�ܔ�7�-Y8N`���Pt���F�=�w%w!�L�K~eY�a��_�J�%���&O�.L�a��{����Z�(�!��h�.�����:Ŕ�۰t�pa�LUc- ����(��[�L���z/��ˡE�|�+���aPc�3#��t_����h`�}����G|����M*��K���ֹ��.�n%�o�] ��Y-$�X���ߵ�]� �],mbo B��������,աtr���j�o=�2�.���C�O������l�##*�b�{=�����u�*�C��+:�^Ֆ���s�5IM�J��!xG��t|����|��*˿ɿ�FZ�j6���M�g��`.�����[��8�{��9l��K-���=�~��yo=W�٘��`{�o��a�jh*�Cݍ	r-���g������3���_��?���m��jV�&�V6� ?K�R���:�xK%���<�G6�oP��-���#��;h��[
z��m]�苻�|]�X�iL�yU�~4M]�k�r��y)� �^�X�%��g c<�äP��n<�2�>)��>������,�]�Wrt��"=���b�h}kh�*k�J�ڑbrN`����˂F,h�����2S�;ࢪ�n��Q��Y����{n9�#�����1��j\E�vbK�C�����7|��{ݨf�5�R͎����>'z?r����H�`��|���!������w��F���qڴFJg��C�SG�r��cJ��XY��f��,�hѶƠB�g/�.ۆ���4@�t�~��r'm��G��*���y��F��� c�L�i��~�F�"t�-΁�_�S.��*�^�|����
��U����R��O��=���hzkϙ���'�s�X@�ڔ/?+c�F
9�K��=E� Xmn�i��&�\|0�˘�5~��V�T���6:��3b�Cg�����.0t������* �ꀀ=�
���%���U͂�{V�l�f41�<i�*�'c��F���_���n=̨����!y!��j�H,G<��n~j$Վ[��c~~��ȵ�7��Yއ^}\�ܦ�}_w�K��,Ln�;�s	f�,�LPB�[�RX{ڦ6���v�oW��Ǐ�D2ihCt6��0l�@��y�z��lq�R�<�x��\ok�vǫ��n�I� Da��u{%��l&�xӘ��r��w�'ۥ���k�rǇUN+��⮐.x:�rLH����ێQ�c�O��� _�5FV�kk�<�k����7x"֋m��(�Tz�fv2]���,v�����K��b�r]/�Z�C�ʥ4����Y5�U#�P
~���E���K�W��,�>hέk�$
^��
����B$D��a�xp����r��*��s�J)��:��,��z?�J�ك�,��ca8p��4��[�����J_�1��3/~�3(��YD�����9A�ǏT��`��Sm���^X�߆�c��v���y\
.)�YA�\�D��)Ҧ��[�y�t�����]u���R�:�%<(�2J��&Œ6�Xk��沼�z��N�Ō���o<Ѹ�J��O��&�`�@��4r,��1@�N1���C4#WD0U���	�l�tě�Q�=�\�:���lZ�|���Dz�V��S�ug	s���L��)	�p9֋�ٿ�g��J���83O�ԥ��>+�s�	� 6O�&�z�Nj<�?`N���y���ACq�l<�1r���ܖ�ʺ[�Tr������3�}3^�!��5�<����Pe�v�$�]�������d�쪓�6z�[��;˰���/���:NM
̝W3ce���}�w�eC��������ki�v��t-?Q�ӥb�;��ZS����)ND�rPm��վV�V�'�J�����Y:�z��܎�Z�Hyܸ�wm�O��9��7I�m\��h.k(�ݽ����]�= z&,��f'e�7+�^cL3����݌ˋE���ԓ�g
�0�nc�{$YD�S�Yo1,����������&޷�FAֽ2L����~e�.YT���q���\�)��=��Z�i������?�r8`���{�d��E���>��]L���FX$�x�MF|��N��
O�f�i�s���WB��Ext�
���.,29�#VN�~��s	�Ez&�C����# 5�
�S��/S�	lQ)����~-B�e�CᏳ����m�-�efn�T���tf���UZt,R����V4�<�Hψ�c4v�/���n:͏�q{�;G$�:�$g�uoҮ����?�=�e����;����Ф�&���=���$��� >���Q�'r��ۤ ���Q�>�y�z������>�sU�~�R��p4�TC�"_& ��-^��9ҌҰ2�;��E�}��A7B��ġ�~C����cI��8t��:!���;�5ԛ��๹i@�ֱd�����F��N�h#�^�m��ը!, ��ӤW}^�]�8�%�0�W��eӄ&�
;�,���]Z�!Ư���|*V�I?����L��{�� �J����:s�qn�)T�
fo�ӎ�%w��L��p��<]Rb� X35S��3�x�]f�]/��� ̱������3?��:��e9OK��kBŬ�b5�H�!��;�i5c}I-�e�.3�h��^:Tg�/�$ ���>뼥?�v'Y�����5�E���w�����F�"�s�b��#�Ĭ)3
^��c>�9�58c�ba��i)�l���d/��)���S�޺�V��X�9���6��\+�ٗ���"�m]��| ]Id�s0�,��.zp���5�`�K	j}�3�b����[8���>6Pe�gpS�_��8�޼���7~�M��K��&e%�U!s��:U��#?�9�#_�C��_<�����*�H%$�VS���3���H�W�Z����.�܈�^�H8<�T�����Bc\�8��mGu)\z'���3b`M�Z�_ȉ�֟ AGc��>E�Ն��q�����yn�_\+p*~��R��^�p���?����]���c]J��$�e��=����w�����T�Ä��h�6TX� ��3�6y�Hb
_}Zگp�Z^���e#�6v��r�6w_)Q����,}�<�3��+�Yj�u#�	��4 � PAr�;�͇�_�ɤ�[�LΡ?����hE��J��7{�1�����{�����ę�W��I��ux	/=�_�_1)!P 4����QTAbSkg�w�/����e�8�5��������V*`y�7��;JN?xK��?q&-��������)���;}{�	�db雌�����8cb�����t �q�F;�5�+$?��Y1}v�]U�����T�,P��:�~��rq�0W\n-5ƩS`�W��t��|0N*ϲ������!:SD��N%�އ6������\�uNڼ�A|L����K���!��Y�p���Bư;K/��-J�w�5+�������,
*&��J@)�v�ә!]o�ap����΢�pzȹ^uNi&�K�X%��s�M�Q�����mj�h�t�Jx�wL�|��������+�9��⁴�@�n<�-��c�i��~|��b�Y�M��uip�����(b���Eg��
����!�b��R�/<��7@��ۏ9l�ū� g6�5,�ʁ�N��^۱��V�ʪ%y�����u���$��g�TɿPA�S?���v��.L��@�i)Z~TF��l��W%�G�P=V^^�q�U��]Q��yX�n�F��s�Ͷ��^�je���΄��
�;�X*�9�w1�����'��Z&ٻ�}ց&g�S�8�16�@���HY .�c!�g����x����&��&�	z$����\ۻ�eHxJ�NZ�PeoY�	�~hS��MpTw�ˆ� �o��<��
`eJmQ��b�|�IE�/ f�,'y�V[1	U�/��� �M�#%�{���7#	�1�k�K\��Ȫv�U���`R�'Gd��V��k�ˀ��L?�f"t���\�>�O>��+�Ų����gn�Pr�n�����DD�;��LH�J6��e(I�����*&3�X$�3�ANW\ؘU2�̶�gR&w�u��w�G�� ҞT���@&�8��9�s�\�;î�N����u4pjA�ѯ ��fR`W`�<ŻO�{�]��Ai�ÍR)zS��(Lq�0��[�n��k�w���7�]���U�l�U����O,�Ԑl��)딿s���Zi>;��]� �Ò{�Hͦ4��6M�د�4���w�8Xͩ��H�6�9��>�G��꣕�A���Ή8 .U,ё������ݶR�*��`A:
z#��Zl"`�����)�1��̿�ui&AQ��l���I"P�����ި�=��|Fb�~�KY�g�"���c0	"LP^����P����<Y:-���w���^�	Z�:F�l�!+X�xL�V[pm��5�ԥ��O(����yk��GV��
}G0�["�P&`���2h�~�{4�vb�6hT�
P*#�̙m˶Fވ��l{+O["��	y�����rx�J[��@X�P&	�BT��,�D�=�{��&K�5E��7E�ov�i{Wd�h|"��2Ǔ�B`,�DBQ����`^�j��1TO�M=^�.�OK�J)l�)�`��8bۓ�ԲĪ� 9T�}m�Τ�ո�=ݶ�^�Y�̉���k�d�>vHoDł��%K{��ȓ`��Kq��ɞK��nJ��q��LJPl�J#i�uߓ���Wx���kP. �������#ܥ8�q{I�]`��%�L
SĄ�@7 GI�:�dq�n�;ߴh��A���%���]��^a5�u���JqS��峜>:�w̾6������HH��I[#�O{���g_fp,�hŋ^w0O�3sE͔[�ć�y#�O�♣�M���?/W���br�[l驘��Uf ���
��]�R.N�3�X��.2��./sꁇ���|�d=�j�vo��^̈��< �2�����+�mf��ɭ��]H��N�݁+�m_�1�"��	��%�1�Vw�[S]-����-_�B�/Q�R"�0�V�`@�Y�Nku�\��ׂ$��S�U�jm��Nܺ�e#;�DV�Ae��cx5	Z�UB�49��� >�8Hzs���p����bki��a}����σ�lEVJ4�������Z���7� ��Qx
��f�$4��_�l��8��I�X�#AA �����7�B���`�Tx܏ۭ��A���./�[�)o���K?�}���:�,���5��X��_�F&>�B�-f�F�
����h�5Gs�p娎�y,w��+aX�'��/.�?�N!O���Ț.[;���{O���8������T�cy-?��$$NRH��p)?�A?�J(����2$WU���_�V �<�����8H߷#��0�hFr��џݮ�W��C~)����8��&ܷ,�\��g������̒�ͻ��h�^��R�:��� (o���3����kd'����y~����^Ѷ�����H����`O�h���h۳a�j�Ѩ��d]x2Z{je�N_ƶ���c��/ȡ���J�����l��F�sʋ.��F �)Z��5	��Z�s6��F±�5�-�|�a����Rݶ��a0�Ѷ5d� X��GC�Y����Ԛ/u���L�¡"	���B�K�2���M��`K|�[�/j�I��y�n%�t�<�����!�&�H���&������sH�W|�{ǟ�GŠ�\�s{{��c�eb~<�r�n�<�壯]҈W
��b:�M[f��,��I�]��� �N�����PT%O��7y}�������@���Z��m�Y��f��i�mw���n�}9 �,	N��ʸ�����,"�����['��Y6]��rW�$�>bo�Y(�(��'��/Kf�S:�D��ih��6e�����H���-@`��޳rEg�<"B�f����!3�C>�6��6S�c2��ďh��o ��m$���e�w|6�0u��a��!s�s{��ā�Yѣ�������7��>ΐ����"̂�z䝻�
�|Ո���%�"S��"h��*����g���7qax�/��k;���3����!Q�yD��w�e�(�GϾ�*�m`R�+�Կ�(�g̤)֪Nj��1/�cO(�cA2-[Ϋ��0�Ƙ���&ǈ���즙��O�Ϧ.b�XE�dj���� ր��*_xiԚH\��T_�����Rk��&�)�T���w8�z�I��i\V�2 �Ty+;|�c�鞄�$�g����E!�zY�:�/����#���ԡ��et���W�v��Y<W���I"��?3���Ϩen��5���N�G�w=)�g"ƻ%_#m��U38�EU�OK�KC�W?��-���c-��/P�M! Q�	��2��0�&�����O�+D)�)%Ͳ�T��]�"Uiq����b�	m��Jr'i8e�����>��#;y<e&NԿT@�J*�SMz���R-ᵅ�6�i茜��"io��TR�Tz�pq����P`[/Ie���X�B��u
`oxt�:���r��qI �.I��/�hg��� L�F���#�d�#Z��,��o 'QP���I��k80N9'3��-�z<p�8u�T��/5_d�M2 ɦ��'~�&�a�۩^�L�����+;���XGh	q"D�q��
"�0�����L8��A��#ky�<=��gز�0c%,B�v������^�|'>�י� �Z� ��y
�� �'�����Hk����$
j���
�+�w�Wv�̩�_���y�I2�ź@U�S���&ታ��
C�wllKk�p�G�Ǹw�9��H�3H�c�*�ǫ]9�)�M��\�|w��� Gh�����U��1Dn���r�jTK��*�;�_
����E�ݤ��v�~���F��S���H�@�`�6>#�Aj�D_���v"���FL3���T������&����AoLL�M��ŧ���$�"�I��
�����+�c��R�&z��?�Gd<dc�@4��!*����$-2_�Z����;�u��s�=Bǩ���u.�i�xRFn
/�7�>��E�mD���a�*�C��8�Z�/��?u7�8c4�*y�+7��(ض�>����@��eÕ��Z�l���_"��,�&�+�fkP�rw�g�-?�oLy�b�kF��W��+�>�Q�1�TK��*�r�@6�欴�%]hΪ�N��qz�`�I�8 �6Z�� \�~���m���r��;��5���	AECx'��ÏB�u�ҟ���D=!����63�-���C ��>�}���㇭�M��8t�����@����S�'}/�%{����wI��h�S޹����V��IAC[��N�Sǃ�z�ld6fG3�Ү"R�Ϫ\��*��.�ō~�V�fܑǬhS��Ĝ�y�ܵQu{�)&uE���%�~�ܯ.�0旄d�]�A��{�˾B�S��5�q���CQ	q�^}<˫�{�r�a��a���19'�v���JD�|Q=ī��ʁU�o ��r��_X[`���Z�]���M# (�r��텸�-�݂T�)/���H��/'�D@w�0�;㷸�M�cY(�h)�\,l�E"��z�˜�ZVA��A�a+�),�J���=�dI��_J(����p�Zq�����YϜJ�]��lK��@<�l�й=>�9XG`w��J�n#o���+%�e�64%M2ξ�@dи9��I����8z:l>SX�IE*
�;\U�OȔ�CF�}��2&uw#H��re��%ι_&��(�g{�>���:}�.��o�X�݌Ed�2d∣r�����lAK?�,�[+�>M�q�|�����g���+ed�a���+�Sm�X�O�Du���$S�+����EL�.$C�P����	:��U��Dx�e����A{X���)4ɔ��^�룃j�3���Fvn���U}HW]a���K_&�\��R�oR0@�N�#�s*/9K����>�1�������A���e��]�|1���6�Z���}|�ƙ���K�Mo@��|Sf*/��8�]���_(�9����^i�n��������=��뺻�)���+�3��Ϣ��I�CX����3�`'NW��Nߔ�� }j�؉�_�~��F9Nb�T����ܯ;��R��w��$�&�?&�=��|�Q�orq��ʠs����?�[A2;���(cl�r��H܌��\c0�:DC�[�lן�g��R!�U���d�	"7���v�������_��8�����E<ᏨZ��F0��͠e�������n�GB2a�.�t���n�F�(��iv� V�1��wgl橯�b�{y�Ni�;/^D{�.�U�@��L�����fH�}��0��
y��_�ȹ��(��*lKS,��,ٮ���"�]�&�F��3"��@�}�6qR:��A�G�'t7rD�^.Y#."�D>\yU)�C�Ah�h ��
�	��NP���Q������2�t��o=�
�B����~f�g�38h�}�1&��W���X-�=F��S�d��ۻX��8�'7_k\Ѭ�I�����U]��lL�w��,��+�j��;52�.&��[�/���Co�]��������Z���L�B���~��<����^�ϡ�0,W[3�Հ��=܋jJy֞B`rM��*U��ë��������5s,��S��`�z��E9Q�mj���� ����(�+����X�s����W���+���J�;SN�|.��q@D֞��l�@�N����:���݆��dy]�\͘�����rE��d�1LFE�ג��F�=���1_;a@�]�L��W�8j��;l�G�t������wQF��$��ݲ=p=9�t��e7��J�/��Ҍ��
륇��ٮ���d��\�+`�]����b��	��y���SW��ůtꋄ>o�hn�jTzЫ�)>�#�jDd�g`'DE5�$
y{^���T�V}!�	Ng�������Dt��O�H{T[-E�g�����D��Oݭ�;�: 灴�,�k8���<ֹ�f*oi�������� ����@�[<�g_ۦ�S(�E:I�4�,3������K �J�z[�4#�mi�����^���,���5�0)G��(�L�\�V��Y��l�d]?f_�W��9���iy�o ����S�Οc6��ZC-+\]��ؗ��и�Y�+�[�ʶ�,�Y��̀�����y ���0�UR�fT7���y\�5�<�qk�7�>�:�'�ed�I7 O�!�)B���rp�a���rG�R�+���U{Y�pA�p#-DjӅ�1H��jM����?e�6q��X(@*����N�pP�a��i�o���#�����/-�`mV��x�/N�Y(�	8��8k`�KM&�L������2J�����S� �iՁ��q ��
���͑�xߊ�[+�����_��B�W�A�v{��A
��Uzb�ã���_�aL�;(~I;�ln&8 T�=����%����s���,b��� �G1q�O���`_Px����"�s���_��g�Ӡmѳ:*���@��W�nM��Q)�����7�����8�	�\�|!�6nA�M9c.�!y�\0!�_�Ԕ�Ϋ�3%eU������"=���ꎘ��G��pc�D�$��w�&?"��B���~�����IV�@���Wg
�����;P�gUsh�ʷn�鱴��)�[�%����I�r����q�Ӥ����lhsѮ��պ�d
7��߃�}#��s`]�����P/�
�3�w{�N��{���׵4���L�ߚf���/D��ʳ3F��(2���1FD+�S� [�0՝�}����cl���H�A�_�4�~#N:�U�҉b��ٙ	n�:�dȫR�&�Y�H�Y��)�����w�K��o��F�g�z]��`�W���Ρ����T�]���6_�VJ*��3V�$\���6Z�	�ǃ�bڷ���|��[|��(.�ٴ�?F�A�����R�pe=5l�R��Yv�,��϶�*g�Zu��b�J8�z\^W�d��Ҙ��f[Xj�w�<xr8�p:�lU�)�"n�D�Gh4�E*)���h(R��a�u��'���^bH��f��&d��6��T8-#�����a�]x,�n��� m�Ne��e�U}s�f��2X�*��\�q��!��l�ݪ�M5�9-qL��W;��*�ҝ��JGv��ր���Mh%W[���`_x��Eiv�F1���������o���f&n��{�g��jS,�ڑ�qP��'�^�vo���f�M�DX�k�
U��� }��\@��<�l;�&f�q��搹/�8�F��w�-��b���Ll�Kv�~?��Z3���AQw��7ê���j:a�_[�1��B�r������P?��c��b.�� ��~�M
���'|�_��3�.C;L_q�?K�VFm��������vWQ&�)��� j+�}xS�P�tO��������-���V�m�4�/��&�i�e�:{,�r�Lh�.�D. �oBh��ǄD�(��M�:���C/�����Rg�#���"U�и__��I�9��ή�p���%�-w�.�����=$d��s���o+ g����v�_S�G��W��33](/����E�lPwB�0ʹ��ˇ~�����)W�g�$�keH�n?��B��m�oq�O�3=���bn#rLF��q�(a�qWp%�uJʀ����?�ڋ�{�L�|��j(Rݸs��W]�@��Gt�Y�peO�K��ja?�>b�MO~����Oɇ~����o�v6D��̋��}�Ѻ�j
�@Ԙ���*�H_�@Ax���cU��|���D�VsmN�,_"F޼����oa��P���g-���*%�Wވ}&��曅�T ���4��Z��\/�!�J�]��(3�Ig��0N���ӳ��{/ ��u+�|�������7	&��nbdUnƠ �-/�O���~����4�iT��)DO$���lB��j=u���z`���; *	-h>�eE�V����d�_At@2>yrZ�@�u��6ÒS^L��P�c�i��)DZ*�*&���L�N>�(�Y]�[H���[�5���g�	[�a��V�!�`E_�o�+��jU����|�|>3��/-<��b%�x�&��E5
:Z��tґ�b�#���� ��� _�3���^�o��}
�@tL���Fm;����w�X��V��X�!	��������J���R���3�ih�(ʷ���E[J]1�A�~�7{h�D\�HC�jP�Vq /*֧�����~Rq��a�cl#��Ρb`�-�r��es�s�������B^��[��_����4���n���U:�ֳ!�V�^ ����Ts*��/�Ą�p@!t<����
w�d�5m�'��G� ���A|��]�I]p��T.B4G.J�Z��1���kmz���	���HZ��Љe"���&}^�J�G�q4�G�J��Y	�,�p�ğ�����38[���=$eQ�����Lßp���%dN	��e��صDI!l�CT��ߞ�����X��M���{�7���6i͹��4�&m�j�k7�zb&� XvQ�~�˗,d��- ;1&Dv��_�o�G�^��m��#b�N����~�i�P�sI�Tf��U�9�T7 EjG�k �3㷄](�M�X�~t��rѺ�\�Z%\µ+5��1��>M���>㺼�o5���p�����v=:����3�K�-�>;;����n.i��r���=Y�7Ow�)���`�z�Ia��IR}H����F@��-��ͻ�X�g��Uত�s[4��X+�7r��{q��u(����ݮT{������#7LGq����nP4�2��.?S��^B�"�Jf&u���}����e�����7];è�LgӇ����{���.`#��(� ,�B�(vn}�)_� o$�H%��b��t.�p$ă�� a����#k�ne)އ�;|���K�:���tȯ��gA��
����T�S<N6�~�RY��dF��Ӷ.P�vu�I����וɢ|�[FA��ļJ�!���������L��/�v���5n��@�;�Y/�����b��X���}�� ��wK-�"[c���bL%:�Γ�A�Jf�uP��s�ﭷ�^��/S>E��������|�B���l�%҇Z?EG��'�e��t���v-�_&��z���N�%�l�X%�ǨF�m��I'2kâ9���j"�˳���`,���∨������MiU����+��n��GD�5)η��?l��c�(TW1x��\f�n:��x�D����O��l�A[�R�ER��5C�r;��E��i&�1��>�3+��0դ��!�o.0A~�~�-�'"Yv䶆^u~������fX^'
�?'
�/�$e�N�$t����U���8=�5Ζ���U��Iu��0����0KG���ءJٮї����Üt1�k�@�?>���=!�v?/%�')�8!\ �E}�ia˗�m͸F�22p��ZXA����^���w��()(K�
�`��]�y��݀N��s!��h#��'E�b��N��D?��w+�Z�"�sj�"b-��>����X��$rO��G�&|�E8� 	rE���Vr_&�>U��8_����i5ߺň�a)�F�L���O]V�w��k�g��mF�����̘ŘPːaƷP<6�&n�n�X���3��$Ǜ<|����)��~�c���}`�F�S	IX"=]cy��E�I�c�	�(�[�V9#P��4� � �
�G�f�Ŏ���;0ur��h�����z�.��Y��+�����{}�����|z$SZH��1�#i
�v��V�˷�T�5�ݼB���r���b�E���!�jH��p���l�;K����jU�"a�3�"���U�X�9�N#}P��#2����G �m�w�TQ$��q�,0W
Z��6H0p��O[�3���I4(Y��,N����/UW�(��iD��O��n���1%�.~L�ұm�A����O�n�����Y�>�,��4F�:�B+=��r���;]}_=%���R�4}��/^�9Ki�$�m���?P
��D��ϸ�!�J�&��	}0!Y�����:{�F�Cl 0��5|qW>�������&���f'c�Z�������h=�$?{;H§��Ԑ��z�Q�����&�����'����xX�ݮ)�lP���2=�s�.h݈��n�,��'�DW|U�	m45PB�=Q�)��-���Ws"�Ab� ��\�~X�"H�;]��
��l}�t\������^er6A��*���l���-���o�*��}ttZŭ�㏷N��;|S�]���!=�+�C�kP��uS�v��"������3K����s�f8U�{��)�\�:��<9�w~�q�1��Ó�=�	�t'��[��170��_ah��j�*rN�z���>�%�si^迶k��uf�'W���$����.�խ0L8v��_uD�![�c6�^�n�2�U}�d�C*��S���}y��	�ص����E2J(���	"�e�Q��(�`�¢�E	?�&TUi繉�u�z����Eٟ�>k���ߘ�Ö�p��z��L�ÿyGK��B��8��]�Ic��p�$��q�s`���+B���Sn&�F:�����m{hZ��vX�1����]���x�[Q�}(�`%�����֮ee�b�<d���l"��oB�@P-UHwa>�0S1&��*%�2��p��~#O��W����ό,�� V�P~x�R��D*J`�"W��s4-$Jm�t�y���pU��tn�6���?�
_R�Wi:-��n��E0�F��?f����ܭ��AL`u�B�w:��K���m �Y�/5�Ju�������L��nt0����+��g��/��R�����u��Q�b�R�rl��B�?%eP헢��A�1v�g.�P�o�m�K�a��V\�{q���K�i�ct���Bd*��&�,v��.
C��A���8��@&�FeN�e�q��� ����;�:]�ϻ[J��Q���*�  �_d�r+�AU���|�����G�8�
�S�X���s=|�����l�C�D��&
��	����W��Q����G���<���C�hH1�Z �*�P惈�I'H��}�W$!�9q�C��AE	� vsq�W�����5�/�K�n�E�3�'�1g�}5Q�^7T�u��K��L��߫n� P�o��T�ձM��;nePQ���������xn��y0�#�l��W8$A�sr�b��C�����$1i��]]�V�\f3�eu,J8]��2�Ep�A:���{49a��[Y�V���;HP������)={]��B��S�ac���Sq�V��/K�DX�IEG�B�!�U�4�5g��2x'b#1�y���B�l�Q級󱁚�]�t��8�Q G�9Ɍ?�t�L<���k�D�Q��S?�Z�5I�Bk0��Lqr�7y�A3���h,Y�x�cC�e'�<��Fm�~&���OA����ȶ�qf�L���#�q����[?�(�--�'�e��U`$�q2p;�,��'��ku�ֲ'��j�u �x����(�6�|ȋ�}�8�#Ma���<���2�|F�-,��&��SKP�h��0�ӊ��6�Z��+���B,0�3��;m�y�@2$�U)����K�b
���b�Yߎ�\'��<�?���v���A��p�򓉗�L�� ���0�/���C.U��D<�# ��Ѝ��j�Ѐ|W�ՆU��Ҥ��Ʈ.\;��E���3��O���T�ow���	7�I�����hG��up�����~���
������Ѱ�D?\�(��� ����<��A~C�t����Y����!��]��]���)\>�5��/��`��ffY�/��K�/�ȼ�xvK��r����ϰ֣n�.�u��/�ml�ƿ����O�gX8�N���ˊ5d��6E	ڣ�j����vћ�m�����
�]Qm �R�����'8�<*Yg���X~�(����}���ԢQJo:(H�����/���ɧҏ'�f�n�W�{׵߮0��~��o7�+ϑ�*�'��#9�\��F��#���(��5#,y�vڋ�!	R��%�c��3���40�C��h���:c���E	�`��Af�d�hŭ��l�-���oSꌏ<]�,3�d�r�U�{fhĨ1�T�IF�C�������W��#���S�c��섔B�>�T��ɚ�&Y�'�c
�16",+�VC��.J�	-����K,�]�\��[m����s�҂��/��x�Л��.Ie�5���1$�����&U�@�G7�_���mr��X?Շ��,D� �chk�i7�Ʉ�lfT�oaw�ꫡ<2 ���q��!������(�y?��o��p$��"����]K6�1��}�'���Q�ϻ,�\M�f���쀇�@�G��kZ�7��P�n��8���Ѕ�o5�����H�ߴ�9^ѳQ�4��@�3��An䏣lZ�TK��j֞2d�����ba��h�J�O��1x��O���(-��4����&[�£��I&�	�]F0��~L4�ć�g�?o�6lk���Q�����@�+�G�(��� l�4+L��]*.�|�m�e���Y���vV�(z~��ع��4��D��ΌBg�v>�+��j��[��H8�ey���s��𒟼����/�>cB(��!�9zX�C�5����u�2Ie�W�#�~q�k�~�_d�~I8���_>����4fCw�f8E=~�p�X����o�ܧ�kH5TOx�E��>�#�)w|qyx+�S�W�b���|i��4�6�Ua���a-W������r���о�=P�l'��b57`�,�L���Ӳ����JDėR����r�POl�}i�����{@��߄���R�g����Q�$ZmO�1rA�n\��_lgRݹ'���m����G6I�	WE��c�9���;v�N��'���_᜗&���&�3�Aס���at�˜���"�V�y'��mr�Z[��D�׹Kr������0j�?�Ӛn�*Ф<Jf?v�0 =��u��ˊ�4|~D�f�%|`��N^�1ff:������cq��d��<�hȘ��i���F�u��pEc3>O�Vh!�$2mr{�N�i�^;ÎyA4�'|#9��� U��X銂x�Z	iܧ��_<���1 �bw��(���<���dZH�8)6�/�Gp���5��
����h�P��d�9����k��Oُp�G9�)sdb>#��h?ߔ*[@5V�:T �.�G�I΀+P����e1�x�P� ��ρ�+JY+Fq��3�cI����K�;��
Q���3�����A�y�>��y�l&���_[l��/���!�'��s���.ؾ�V	=Ixڦ��܍�B9pa��9��t����MVR;�< U�X�#��ht�~����h]=짱[I��u�Q�KY�}3��N��#,�r�h�$N���F�;��}�kBn��-��P�>��_��ⵙ��ѹ��&k�f2%�e˽&Y��Tw�7�,I?���Ձ����D�~�5�c4 �>��o�{���w
�W�'���T��v��|��a����&�=<˰uN�辽���WO���Pj����	�:�t���s�8I��l��t���Peùt��D�%ex2'^��8=ٹa��ݵV���0��~�8���"��e�S(�}����?�x�y@4�t�&�C��K��2�_��3�yN}=1�°�w��w�������w`���s\,u�K$�76�	��J2��q��*��o��FF/ۼm��=���~��ʈR�,���b�-ͺ�Q.�-0�)�۸>�3K�ږ:�c���|�x�Kv�_Ggm��9]Ayu_��b���B���Ns��gp�8���c�6�n*ڵ�ղ'J/Aj��˼ȧ�.ٺƿ3�[[��x�B�[��M����N��e!a_�4��[��#�%�R�;���;���Az�_`!c�z;�7Ub���\[��%���*�)��}�m�(.��~Ox���I��>O~6׋��{ꖡ������h�s���Wq��[4,���d�X[i����1E����qpd��h�:	��8�4�j&y��Y=����|�����L�z��]��m���+I.�ʡH-ʦ��x_�v8�7t��]�M^�GH�J9�����23��e��u��,ӥ��������8�uyh;&PQQȸ�OL���N�qc>�\vU�ڧ�R?���T>����<��/���-ThO�Y���<UY>�����A��3���"eG]�F��H�x�`�'��\=��8�C�GSo��S"���T��A��v4�cvQ�J��Ըl!X����M�P��|�-���͟_�L���tE�FT���tc*R���밗������: ���ɳ����3�N�/վ#��l�N�W� �`B~i`�r�{c��&���O�� %����"�;�-��4����]����DEj��ap�^bUT�*���Y���.��b���Ð��j�璀u�&݈�f�lt˽���Z=�uNc����]�c,qeW��6
#~���ʑm.���]��P����昁�Z�2K�U.j�EiD�����"2,� ��/^�!v�WLf��P_�GC�8ȟ�(i+ď>�]V&�̘��\J� ����k���:�Q>sA:��А�Wԑ���i�� ��-�m#'��<0�3��[k3��4�v��>;�6�F�j�GK�%t�A�,Z#OUq��v9�`0��1@����v�9-������4��Xv��4��-�BcS��C��?��0@q��,���G;DaAl�q�ߦ�ʟv:s��
h�ܨ�θR ȇ���2{�7���4˽�,�_�t���A��c�b�߆�76��:a	�2t������A��~�L��;� '��_�J7n�B|,�0�t�����|��?��<�AS�7?Q ��7	���w��P�K>�
�^KH�qS�sY��Y:q�6��q��[ݛH���*s ��J]E���^G��}�������f����E���Xͷ4dZQG%\��l?��]4f(�x��Ӆ�k� ��Q�!S�C]gl$lOy�߳Z����"��[�#r����z��!2;䲎����<m*�W���c2h�}�0�%�cx)�9%I�S�4���m��:��o�Щ��).<�'2��I L��~����}@�7HE��	k_�(PN.�98���s�]!wb�.u�s�.1�}"'/�Z���i�i̓q)8�.w�e���I����)=D�G��Pl �I
{7���2S@��.^��j����{���?�Mg�H0j�iGZ�DL*\u���''LNF_
���%;/:A^!|��Ľ��;��"�W3=f�j�W��V�tZ��,B�՗��it�~�#�K��p���Ơ�Y�>���&��=�[J9J�2�C2��F0�դ0��[55 ����+�m �� T{h�y܀��(�|�(y��T�{̋�X�Dp��ܘ�����F��S�8q�f���_BSY��np��pt-�k�g����UtQ���� zJ�]����V�`Cu. �� �E�;m���n�fY���w�����<~N��;�aQT:���2����~�yJ*�L��J?���NL�l�lF��|PV����?S�
"�]_c~p��(�쥨"��UP�T��b+xC�4��X�\(�Q8��<N9u������J�k�k��n26j*KQ6��B���.Шr��Х����Dv�Xģl%�u��ک^�����t�2�^d���h�`ö{H��������8�'oH	&�wzX��_�c���O"�1�o.�D	.��A3�_���j���P�	�_�|�|�)����G�E�iZ�u1���f¡\������2��P�7�q�AG�œVK�4��^�Y��k8*�Ѣ3����a<l�|�,/���;L��.g�	p̺�h01jW��S�c�c�;�#AR��`�_k��vƧ��g����5�_��ƈ����
Duru(4�D����y��#���?8��qV�ِJ �SΝ�g��g��`�;a�n�_�zI�k+�Yf�^?���� q�<f���l��W�%iR�8�E��>eI���0��°\"�GU���t�Wg��/+7#���|q���M��Va(���K.7,�O��G�X)�B�~�o�X������̠lu��8�� 
�X����+啶�������V�嗝z��ƴaY����+��ۖoǑ�S��ӫ�c,�\)��gC���M�iؓ�"���6�IEԔ�1��K�pL3���u���Z0^��K60��9�y�[�\+���Ai��C;�l�⦻�#��F��S~�
_;�z�ߗ6A��EoUCo-�3�kp�1���Ӆc�$o�M�	�� �������P��ke�Yc�#������T�G	` Cı�؀Tk �!�`--���T�'�:^%�܋�X�'���s,ܐ�H�jʑ��[���~tI/��V����%0D�p�U�v�%0�H��,xE��g��`��4�W$�VޯN���=�Mй�-��&rA8R�YQRS`�`�O]ʝ1M6e�L ׁ;
���C�<
b��b&Kw��Y�����}w7�z�?怼*ж�w��D�� �[_���Q_8�P�#������� \�y>�O��@V	@�I!,��%삡"gV"u�jް������*z�%��.�-�{����$f��#Ύ�m�}t�?�O���:ʯg�G3[j�e��� �&�_�6��
��aτ�L�'���I٪��bP�MZ���Ҡ���XÔ�����$�.D�#�Q2i��i|���,���b�nTV�^#��Y<��\]�+�w�#�0��ma1��k[��{�4���zJ��J���z�W�b��*�L����!-��T��J6�g�\ɶ/�t�	�O"����˄�����rCQ[���'����Ѽ��:$�-KWP�e7�_���u��/��P��&�>edԺ9	!Ol�my���ğ⏈��X��� �y��L�Z^nU��t�9b�ÖuV�-���~���s��K���d=߰l��}���W)#d9}���A�ƣ{c��� ���f8���%V�:A1N>jO�d]
�燅T�pT�����:��'�70��u܆P�J^,�bh��毁"��������+���t6Z3C���]#ũ��Д�i�G-Szo�N��'I�5����Ea��1"����S+[������k�ÖD ���t��A֌�UԽ}ё��o�ԁ ����;4~��5j���X�ߋ��S�B����C���{������a�
�p�*?��<�΢�������c�X�j�6]&h�JDp���r+$�T~����j�l[��
[�~о'
�xh����r�a�%k��tmJI3� [��ڽ�|�9-�]��KT��,�SS%K��dLw����@%���n�U�K�s�9I��9�7Z<?e�@wp�_u'�(� �ԧ�d�1s,`~S0�T)���qa�>��`��hT49NN�q)0Xt.yp�]����(���<��uI���\��o#��*o���Ѣ:%�1�D�%��?��{��^��Q�����J>ߚ�<OUs"�H���B8&��o�Nsj`�h=߹ܻ� � ���^q��+Χ�"���(ю_��Mby�zt���{u�������>�:����A�;ED	�ݬf���yK�*��W�2N5|���~Q��Q'щ��.f����:��{6�	T�{��;F�8ڤ���k�o���r�����A��5��ҕvs�>T[�^���]���8�D��o8��4U�ժ큉z;SS��O��GJ��u�K
<Ц��b��U�iVo��'!��M��BV��0�t�X�0�3O�<�p�f�HT��@DG�,�?JPR��>J��'�V�/h_R�B0 �P��&�������TT�kuֿq�R�����H�ۢ�=���s�L�'��nD`��%n��y�� �� @�ܱ�����^M6��C\q������eyB�%T��e�+9@�Pw��{��q����Q,��Fx�ŗW�������)�9FLԷt��-ܤ��`��-^�y����Kb���̉RH=���.(�*��3����ut�W���TL{�<�3����rݰ�!,iy�Y|������y�����Z$���,�-��b��ꭚY��).Du���f=  ��3�C���ˬ�	6��yŤt�����S�	��E;��w/��r�Z�/;��3�=A�f�6�I�UXU�{�8+�+�Tv��#���}�&��ww�i�˭��j��r�L�d�Y��f�;l�%��2��9gJ��A~%�3]t�Ǡ�������;���c�t�؟��b��}���դ���@�"��Ԍ���$V*��p�;�W=�:*�����&�س1�M���i�_�q��Z��q�4�%5�>]�b�j�?��*��#�>�`���Rٖ`�en��4���)�p��^�2�;>���{���ޞ�un�<��w
Y�\ ���"�
<���I�k��Lp]['��/FN�	rU�vԞ�b��6�����	���t!�2�!���{��|�WI�[��`���:�]�@M�+�5-!����kAᔠ���o�A��C��W�+����9�VJ����lw"⢣�t��G����/t�L���qA@����hZ��L��0(��ݔ�d�_!p骞wI��d���|r���L�����@�Ŕi�֬8$mj�BU��^q\a4��p�!{��K�2�ygNܙ���}n��"�K4��f���Y+�ㄡ�����HjL)�GZm({�f�OE�zu+��i�Z�dˬz)��ʊ�4����g_� U� �D��W�Vþ!A@��%�^��ձ���կQ����;mk�>Qu�!T�2f�Fz>�v�6ѿGxL�61���㳰`����%k!��5��J��f�b��r�%uc�z��n/�XX@�Z&/us�(g��v�_�"���$��Ð��%* ��4�II2Yɜ_`�i�5v<i�0V$�u5$u�v��V�*�58�MUf�?G��'˶�df� ���/2M_����B]Xwտ��j�.g��k�Ͱ�Ds6fb�Z<��$(���0ɞ)�ܾ�.$p#��؋Z�ޘ$�MY�E��&$;�����9l��Y�<?���������] �V�0�7X=�)�q����p��{+���u߱
���I��ޔ]
��0��bSlYF��� )�eUl��X�]B�c��'{������`����p�U��_Z����Fv"��s���G羦��}]�~���O����'�g֏>E���R�S걿���iO�}����5wx��s�Vx���(�"SW5.��GP�1�2�a7�gb,��޴��c0:�:Ҭ6�̮���Ϡ�0^���G���F�MM����f
���ê3�f�I,��"]n!dVԲC-Z| �X)��<+�o:֭	�^��������SׁI�+�)�����3��N
@�se��o�5�bm*�j��UQ����v� M�6�hz.���(�(��M��)0k@��O%���!��[�_X��L�@��=r)�FMZL�<8��{������eћ�jQ���@��tlKS$����e#<|�chW���c�¿F��~�Gf`R�e@�ެnv,���IY�	�Y�	�=�S����<��sy�LZ����*�zj0�D�!%�ꅀWs��oc���vB�gQB	&k�܉����/SUcU{����]�Z�.�� ��\\/'RY��,�/���,>%�LbT)~ٰYE��9xbk��>T-MY*|$�6B���z|s�W�C/��oƿ��[�C^���7��tg ��&)�!q�aSS��4?�ix(X c�*����j��I�����]+�]�nؾ��ĳw<0ټ���#��K1D�����SC���Z)� �\^�0�g�"c�ļ�3�<��q(w���� pV���$�h+z)�ء�k�����IT��=r�Q�3��8�D*�f��k�D�9~��i�� �,�D53��0���ŉiu�q�Yݝ�Z:'������#�0L�p�Uډ�}~����5�"yL�3�|��= N�u/��W��F0��Y����u�X�z�EG4u���������uxM�iqp�Ӫh�)b��B �*��L;�a�m��a(�V�d7�V�ŷK4�9����2�W%<6.�lvȉ��,=�-�j��s�uMꥌ+�r~/߄MX��>	!����dҟ�0K\���Jc��mJYXR�~���'�Sƹ�K��_�@IKv��=p�s�qs���Er+��&CI�9������)�lT�z��Ҩo0
�q��'sϜ�IN��V��Ǝc��i�O���<z����uI���% �=��A��A:�DxU_@�k�/�J��5���i����,����}\`�e/9k�3W֨�v�l��A�sy�.Z=�WZ�� �J�au �s��(�����H������� �Mi�q� *�=��d�we{��U6�^�3���@��T�uhm%I�������t��ޭ~�g����Q{��.C޽�gO"���%i���c���4�P�W��:����"*Cly� s;"��W��	)d�}���/������
y�]�[��<���-��t���i����y�^���n�Ǎ��VY��-%��q1q��H�!s{�mR� (�b���_��yC߂/�1\@ K�K`P�����Y����Q�~)�=�-�k������c��f���P}3���i�cS����@u�Ӱ�C�932֌<�z�"���x����3X�)��\���^J������}���Kn���,+���h�$C��:ʚ�Aenq�$���f�)�S	�"�es�j���'�%^�O���֥S$?FYJ$o��+rh8;��i?��W�QmWvr~�)ꅩ�`�)��O�rsd���"0�f��7[��s	dV�*C���|oIaX[�����N�V-,�~j� ���7�CT�U��9��g�o�Ն�·���4E( CWմ^ �+�Ж��Ɯϰ�����!��Q�l�5���O���u`dZ	�%ﵗV��(�ʚ�+f�Sb"/�D���PV�}�x�[��,SɌar�-Z�>Y�;�&
*cd��:�ݧ{T��'L�y�;]��a/�y��識�9�xR��o��O�`xj�yK�#fj@y+���Np7Aoixx� ����i��$p�ʨO*GO���������3��DoT��C�2��0^~d�.�W�C�Q�9�!����[i��l��Ź�S���*�"� :��؋�3��C흿*�Qs!%�ߐ�h���mn1�Nҿ��/�c���a0��p9�i\���ǡ��}�u�b��^�r������薮�����=��JS�O�<�|�k��x���/���5�W,SaL���>y������!���{&OwW�)dpd��r������wc��lM�s��Lt����L��Ʀ�Z�X]\�H�� �i��"	)��g9�P�.+Ü�}pii]M1S	��M���Y�F;��tV�9�M��c�������Dߞ���}�b�h�,�����MZ߁B!����B$�! ��܄� ;G'4E�0��#��#���%�ϙq7�A��q�ħ�(�V	�{�E�H ?y�����*�$���A�A�\xt֕���?���,�j~R�q���V�a����J�'�ec_�us6צU�M�I ���٫:RA�z�?ɖ��k+�����#V�ˑ�Դ,����1u�W�������ߞ�����_-z3D����A�~a�V$;Bf�z I��P��Jd�����_�$�a=��t:�6��N�C�Vt�B/ ��5��^\�hd�� ���x֎�p�}���&$�q}�ڷ�쿑��������lEa�=WXK���4u���$r���pu�J(�(AÜ��Ϊ��Ų� �ښ���4opmb*�3T�iFo��������0{�Z���m��YD�	��lV�������3��1EL�t��q0R���-p����/�WSs����S��ã+"�<x/����T=��c��m��`����6Ct}r�SBƾ��+c�br��_���(#h�����w�W۪�di�xq�r��m��9��)��p�Q���ݎ�M����A���$���6.��tͰ�8>��7���6�jb}}�P"�N�|�v�IP��F8,�'~���))P��M9�;cp'��Ґ�;Dqݮb�O�5�2a�K��!���|�J2�jJ��;9M�)I�{�r{�L�$�L�񺺆�%�^L�� a�{i��(JL�q͏�'u�Wn��_-x(Q,��m���Dl��!nޮІ�����%����*���܀�e^VHK��_���1o:VO�c�� �Tյa���=9�V!)*�f��?�w'Y8#yxyd-GMN���W��׷�NړE�e�Vߠ��:g�&��vB.ߌ-Uɥ����n��o��u���)�w��	ƃ����J�{xD�&�G��-��e��2�>E�>���3\�('u�M�o'�Nu[w�#�����̇��o��93@��������;;6�\A�z� &+��v-%�)�N�R_�|�ިy��a�Ds����E8��[�kF �b���U�W�:ҚP*��)�eM��"d��;ǭP�Ҷ.#&�P��(AvB^���[��{	w���?�ޗ^�P)����b�"6�j�����Sx�3I�2�3ķ�d���C���x�N�SnT�<ޕ�
h`j,�0 �F�v��ͪ&�<W�Kn��zK�-�J�>�}����ի���ɠ���g������x|�`�b�=����B��q}���{'	XFw��M�r�t��3�c��a�7��?��ņ�^(D�sdM|1{�t0��������>[;��D=�kN6��d^o��g%�L��I��Ё���A�@���-)LmOe���կ�:{P�º�����zx�8�X6j�w'��������r�����~��__�'���l\���*����ux�O׾�L(���1�R�j��E�!\������'�>���B���(�!b�e������<U�a��#"�SE���y���@�:f��q�����2��ү�z��PHF�M�M������E
j��8������0qq)	o�Ӄ6$��%��2Q_|�C� ��K���̑�mm�U�{z����aW�O���iߚb�Am[~����a�+p�>��і�#)�Z���nX�*;
���8�����2l���>�%��j����S��!��p�f�9�й�&��y=�^#fo���7�[���c�ڡ�	@QI���:���xC�A4�V��(K:'�{@�J���\(4�G���H��Wyd��J67�(�m��n�)H�f��������ڷ\d_�H9�T>��Y�s��`]�e�U�SIg#0p��6@���7�%i��;GT�^��=b�嘗��>��g�]2�Xdk��z�VuY��R9f�����c��Ab>�^��a��*#1S�>������A�3$���<1�2e^���<����F� 3�^�5�]k&<��۞��b�Z�8��T�,Z��-Jm8@%h��Z����~.i4��_f��m?��J��67���C��^� �!��`wJj���ȷ�xk�疴��襫�vl?�br�f���~D���ng��V�'u�S��v� 8�m��t�s��VE�^�,�;��5��zQ���U�p��qPs��$���P��U������k����Ӧ9����T{�j�Z^%��#\�Ě������:`n��V�{ ��uB��pA}+����7t��� �<�p��n��(�HY@�T�z��b׭�f`И�~��[�_e�2���?�o�1an�����E��^�>�����y0� =���Q�Ӭ�q��ƢRI�Ɯܢb����b6����w�n�Avhs/"�=����y�����@'/���ʞL>�ڡ\Ϗ���/:;�җ���W�� �G�V���5�;e���5Ё��3�x��Txb�?�����~��|�����9�
X$�dBW��ᥡЬ�W�pU��@�ŧ�9x�X.��N}�N�7��ubA�8 ^ �;�t�M'�����%�@Ē3�U������83fam*b{A�x�+m����$p}?[S�>3��T/��lj>>S'GNٛ��{�9�K$�{K���4��ɾ˥�؏E�Yt��E��rkR�	/�m�oiј�G�cF�#z�D��!r
��ys� /X%�Cv���?���ܺhn�I/A�[�T.`�86��s�V�uT�E5׶F��#U�����@h�����J��Ƴ�_�a}Tw��ߛ�I\5�Ո��1���	�Xb�/:]!X�cɵ�G�����c� ���Y�&m�:qˤ�o�
�+������.D�����i^��ҷ�t�Ĵ���(TL��\�y��?�!��{�qTQ�t��4�#	�b9=s�� *0M�:�"������o��o�SG�T������"�q{b�>�����ԧ<Tf,�;=@7�5PYx��\� �=��K��S���bh+M�/��A�x��}ʷ���g�m�[K%PmG1MGs�2��@�������D�5e�o����LY��7A�I�<�%�����TQY��Lv�OL �4F�:���rѧ�E �Z�-wK<@�xEc2]U:p�5��n�s�lx���P�ܕ����	�p�;���`b� �s�M��C_����m����K�e2��}@�]�v�f�٣�yhP�(1u$$0N��i���L��&��H��g��I$�H������������zN��p1����n�2%w��Z�f�o����$iE�Ԉ�D�$�8�: f���|rw�	���f����?X�wzZ�^�ސ���4���zW�8�x]�A���L�U��k+��г`avWN�_u�N:�۝}����{�2���DPœ���^�ģK�3�lV2���������w�k��	�1���{(-�.�쑧Յ���,������$͜x�������˨>�W��Ry{$��љ�}޽���ș̓�T��>�w;�yl����TI������l��e�#w�D���y�;�%�Z��������+����A��՜�/V"'��T��9��;�p��w.�?PU�L%��;�r/��V��aԇ?����wv������y��;�������S��z�V���1hx�{��g�b��Q���z��g!�C�o������A�~���]��������'�A�M�Y�{q�s�ʹ�`~�������mS�-]� L4��8�yJ����@M��Ϥ����K6)��w���T�9��Qto����Tå�R���ܗ>�}�Ôt}��i�f�:G�IsR�LA\ɷ�#��'K��S�0ja[(�޲�ob"�BS_H�N�����W�����;!$�tH�;-��AwٰhL]3��o���+s��=|�횓��>�U�"��� ؀c�8�s�����c�}L�$g2:JS�i`�ĖG�j��7�9E�(2�����Z��
�rk]A��6�-x%�	�C���,�;\���#�c��>�<z���n�)��2׊߉�~<g���f+yg�8����%'�4��BoyS�ޑv��-�n=�9���M�S�,�<�% ����Rk{\Ӭ(�f��i���i,��4��r�V�	�����U�&OVE�D�vQ�V�$O
�1�.�h�Ǜ��(�:ͻ�I�I� S�{~?>��;~�4����U1-����4|���m�	��iP=٬���<���΍|����<{� �+��ŕ��Y���>*>�mSy�ݘ����#F��'A5#\Q��Ѯ��mS�	w�zH^KR��D��?�sj�3g�(f���ba(Ө�ky[.��=��#�|D>%��孂DS�SM�ʣ�k�y�`�Q�ht�լ�h���1@��з�g�\>��&�������K(�Si߁$��T���ki��~��iqbT��P'�ҳ"��¥�����%�rŃ�mcp��۴r��[g�Z(/��d�ߴ��!�����z�9��|i�b�M��\��c��n��օg�k�Z����7��ʊP"S	V�+��>�G������$� ��b�`C!�	x"7��1%�p"�g�gz�L��;�9=8YN�aZN5�b*���m���H�v�%n�nv靝q���-�U��,�BM���bɢ��ɔ�Y�e�y �P��d�k4c����:�z1#��N���n����y�ΰ^EV��� ��)����j�5O���1�nIk�g[yS���5�����1��O��:�Xd��S��	�ZIܱ�_[��h���V� �T�'�`�)$�۶�����>a��1u�e1�__䨿t/f�]l�.$��Q���F�n�jߡ�eG�����)V��i1.��n=�����Ϣr���r�O楝���(
Ţ���?�W�����[�¾���)M����4�`M
�#�����'�>�����C2��3ăށ�?.�k�noi)�j~�y���k��#�^nKn���B�(4�5�gXt���7�����,܈xd��%� [s|.�G�
�%����hQo���>�'V^.�7���r`b&NK��5�v��7�uP�23۲ţ���P�XOE�ع���/bOt��o�����(���_41�E���=�i�ή��O=���
��̔s ��kV��6�|4�L�qq�=T7>4���>���\q����]�th�B��5A�u��8���ԶV�����������	Bg[E�_e��a8V(��nFl3M�fu�eA�,�.��Kk|d�\�t
}�C9��4T|�n�lQyp�ݐŷI*�!��S�=G�hmCc�u�zw��ά"S�b�Z�a���Z�aC� ]�ߴ���Gj�pS�:25��yl|�v�u^��u���:ۂE�E��|VN�h�dlB��H%#�R`�
�|�Q��[�� �w+�d t��BT
T��@�X���wr������֯J�V8:/?����T#��6����M�� �bj�a+�P��k�FrX;�C�w4�
�d��$�._�3�u�%ەR5 �k|ўN�>)���D=p6x�~��I��7O�"\�~lg������j�݃��n3y��n�TZ��ZS�'z�:Y8�Z0Ź��'��8`м8�L$�+���U�24�������}��P��6B���H�
*����Tb���o&�2=��a�c�MU�MIq��@sD�t�oznl��c#r� ����9@�&�Tc�I=�&�il��FZ�G�6A���Ou8	�nu�]�<`���)�F�%!Z�r�oQ�u�Uhr4|�o�Ԏ��y9���ȉ���F����B�$�+k�;��C;h>�`��ܳ�l0z�!�.%�=�HI
�<�ƙ���cI(�eґb�$�n��jCR7X�:� �&3�\_��wH��T�mҫ����9U�-��,3��K~�}�2��C(P�)X��
 8���c���+�8}��0d�����������+��7+�p7b�}܂7�����T?Ma����G��"���cݔ���c�Ra~�S)�ć��_F��g��w�Dј(�I�{e�:}�޷�A_�3oX%j�(x��P�q���R�Yz��=�ՕZ���m� c�G��� ���O޳�F'ʳQO���� �?��ͬt��2BقHupC&��ᮍ�"�������߆�����W���J����P/:bU�1�����,���R~����,���d1�����#����l�d�'ِO�V��Ɓe�N���6����1�������ǈ�W�_aTt*x[̘R����_AU��y+Q��.�O5G�6���R����ep�{��w ����^[Έ�7�Hl��tۘ�sj�q;~l)����S/H��.��p��W+ɔ�?��FC�+��� �(��qyq���\w�w��8]4�����9+�9<ϩ.A�s���&�sTsSa�@�T(T����3���9��)�UH���k426K��2ҿ������!�Ҟ���-���3�	r���h�؉+��(�Wz�vG*-'���w�ӗ�����LyG�Yb��9�Sʹu3�{�B����A�#-Q+�k-N�0fY�ѽLyAn���5�Dc�?	�{>�k�aU��\�y��+�r�|;� j٣��ʶ� �'��n��ٹvef�@�?T�s�����c^%DF�kc��iD���wƖ
����&I���%-0�H���k�o,����3���Ȩm�GQ�sz�����@�}(n���=�*�8}�+C�⋏�=/�"����� �pG,'�7*Q'K�9�۠�����~�	��p >*��CE*щT:ԧ��\��ߛo�Q5���C��2I�X� ��4�nk.���1@Z�9���	�+�~?๣9�����b��?��X��5��,��@Gd���IA*#ߺ��kkq#'\�wy�,B��`6,�����}�����6�T�O&��*]C����:q���G$O��M"j\#���|U�=��vԟ�5Z�������� �S�:��(v���>��F��GސoO�Z/~"�L��ʥ}�#;�I�e/�׾�$��q��&�Q��R��;OM�G��0�h^b�ɫ�+�2��X3f�L���I�!>�?nd֛{�z�[�X�<�ûp8g�;�
2#"k���ec�0]�������0[�)mH�
���s�nϐ֢�?�g�����)����1ۑ���=����$A�夠�WA9�C�V���{<�~e�ƈt�/x�}vO@��^O�����)�<�<SJ�#�����v	�W?�X���>K���>��Ӵ�����\o����߇B��a��[��= ��b��p`$���g<���)�'������H�I��l�t�1�i�t�/��@�i>�����U&�R��T���l�Q�@,ŝD4nÌ�4� ���h��&�G�f��D�Gnzȩ0��(GN��<*��h�o���;,ad��-��.CZ��?�&
h��rA�`;�ȭ��})L9.tE���Ѕ�n��2�� �:�K"�u,���j]��e��`�	�l	�,�����$�.���+�+h�����ا��	���ڭ(_�&�Ⱥ�q\�Faq?ݗ���� ~D1 ]·[m�Í�<k�����n�q{%df�
N�FmsHڲ/�m_[;ŁҸ_�N�i�p��`Wg���NX���A����<���k����D2��;�`Hga���W�A�b�-x�,/Z!��������9��9�k�(P��=d����?��Y�-2��c�V i�)L��^�o��ϦC8b�r���?�Vrhг/��2��7�!m@�s�C�Fxf*�!��\Š]���3���Y>F������vm">hY��H-ߟF2,�1�����=���TyF�����G훕(�K҂[��{Zs�)�&�M�Y&A�]��S-*�L!�0��F���P3h��tQ�=��]�x��}D�Y�T偁Ͻ�R��T��^r~5.+RѿD�VιW@{�W�����X��8����d�3/�8�Qb��Oʝ�e�6<I�?��u�����Yd��$�)��Pm��d�Kp�v` _�i:f]F{F%�.�!B+�|B�5q~��j��r�E*�8�#��xm��2�_i<�X	D�O&���$��bل-�L�h�HB�1\Ĉ�g���KN$ �<�����zw�K�*wW��D��[Jm���[l&ʌ����K�>1ш�y��5}�e�K�`�H����Xsp�ѝYV�)�"���1�������nc��	����V�u�D�1,�2��}4s���8�����K��H���#�ǆU��vîj;ͬ<�cO2�War�j���OFL�
yM�!����{r�j yB�S;L�)��*��b�����aL�E?4!&(�����Y��w<�p$��-n��F�`.�^��m�z�&��a_~5�+��!f�o�'G9��5���w-���^�ayX� guC�8�"�(�7_u��/��|�Q��fX��嚙Gh�I8�s4�q$Hu�7
;
�,�U��*�»���3u�������4=꟰˦9���T)�q�q��.�BY[B,�~��(�>�VGH�~g,K�
��И`Kt��h�9�g��t�އѰ�|iw[{�z�H\��-	���+��ȂAa�@�\�w�fmE1����/�q���2�J���o
����cE�
�ab�*�����I�1;?~R�"��X�u�0"���T v�o���ER��lߏ�҅z����#WJ�� ���3T9J�<��E,8)��l��_D�^�'p�WgG�U&�k �ULm*�8�Z�~N1a��� ���"$��	�(�{�DYY�<�du�)��d���r��v�q�UW��m�l��t�Tۅ/����[M9�(^תi�g_Q��\��<�Y��6�j�tO[ɢ������@��g����,��۠ڵ)A���+ԥ�g.=�DH��s%����w�Q���+�;��o�}	9���ͮ&�*�ho(��M�ļ�[�HG�+���rx|.�|�fQ���њ&]]5Kd^#�)�q���pG�r0-g���C���0���P�����X��,0DQ1`���������QxA�Ca�������,�	.����*��߳y��0��=�~� ����T���IQ��Iy�VGȶ���>!��E����G��)7^2�&�#��oٵ�r
�ӆ��)^h2?��˾�ɡ ��p�am.�~����,��j��s��KW<�F�6-���(�-1HPit��Գo�Ư&�S�q�c������Ǆ<�����:��/%��{@�t�N��T4a��O������G�J&��/p�k��U��������n�_30%G��o���_|��z�B��1l­o�^��RG��� <��@nx�ZN�<w��� SB�0�nA��bx
<�K� �֊:袒]��φ��:�1��*�>:�?�`?�ⓕ��i%�q�l'�z�f1۩���A7���u3���Qb��K�Imc�z0�a=F�\,5�#z���4�Q��T�C@o��'X7Ke7i$tw�~'~"���$�J0��)KmH�,�Y<x�	�V̋����1��0�R��ȑs����N���&ߩLD*h����t�\(ʞ����E>ʙ�R�N��U�H����ͦ�H�/FL�g}�Wm#6]k�a}�y)�cV��?��j�P4���{���+�X��<�����P.��,����� ĭ(���;h�o��G�3������]�	��t�݇�Nę �ޒ�Do͞���z��%m%��=���Rdf&o)���tPu�t�>�!t�Ȥ��>���T�\�7��1)p2� �϶��Vg��r�$�M�ȑ����u �T��ې����Z������3��v�h�d�R���:�`e�5O�m���j�bq	�$�6O�HeQy��g�8n�s��N����+xa���7����ʹ�\��)<gw�y�� �o��
Q~''��ܧբ��o��}+\�:�cD��A,��˃˭�,���\c�1R�?9�J����S5����1�K�cD����E!h]s���֧1��Q@�l��l����ϲ�p��'82��F�xkx�˨��y2���W�1@���.��R. �	,�D��?�?�񵡯Y܁#��'�vdi���u\ܭ��P��N�j�ܴ'�N|����+�N�s��5��M�_�Z�#7r�n�<�)���
g�̾%�ߐp ������ %웅H1�f2n���6g\ג��=@�(������Q����G�ƾ@n�c��>�J��߯4)���	B�f_��~�g�B3�@0�`P�y�A�$��bŐp�U�-�=��*����6dYXa��>6�F����4>�>�M��n5:nNӹ5���R1����L��~D�/�`�NSZ�i\��na�Z�H��C<��,'Gt����R��i�>�t���mm�~�ދ��~��&�^���
�x�q�\�w$T���9���x/2����{~���[�mm�E��
��5��~(�tg�O0������tgH8.T����ݖ	�Eh�2 �|&���ȁ��$L�m�E�
�CR�m�o�3��l��:\���_�}ϟ��� ���+�d�m��*�-xJ^~욏��foۂ��fJLR�=�Xݻ���u���%�oH~�_����6��U������i�<gz�b�tG�L��W&��7�w���v�K]�����؎���CZ�5����d�>�ˮ@�{T��"�7���B�b�KQU��ҞH1�Ʊ�~@q��Z~'�OVvʱ<���_��>��X[U#֊	�0����w�Q�r��H6��0���Wʂ�����m���l�c'[��(��p��Qό
�b�#i�$�R�l�㎥��I�)(�2
�V��0$A$U�B0�j�w�2l�����[��Oz{I��И�(��LN5`�x�qho��l�6��F���@u��`��~J�=�7 �h��nLx��9�����ׂߟʏ(:5���P�o8+�`6�Q�X8>V�c蓀���B$�ʮ�7hnL�5j ��)�#b�ey��bO>2~���l3lh��GBc�uRN�f�H5 mP9�i=��c__�	aϟ8.����������}ު����'�um�y�W�!��~�kf�#x%����82���]o���m��i��|�q�4���6�7�
���ܲ��H����?���L�i4k��|� �;�a����4�Y&23��xNT�>K]�K'�=�����O6Y�����~�x���	�ѵ������f�M
9�CTlQ�� �D-�X�	�V0�|(?y��?��%��o�e�>9e�=�`t���נB�R�-�i�z>I��Xڵ��G3� b�[eg�����������a�Z�9(g��_��Dߎ���w��}��i~��
��MF��jY%�3��At���Rߩo�UV4����_"MZ#q^{o��}���(��n9�i�&���Y|qN����/]�x��B{����.ǘ��G�&"=	�D��Gox��k��7b����W��ػ� ����]Q�^[�B��3����3nc�GGa,7�o�vw/OM7��5��"ىkzo��T9�X�Z�p�'޵̈q��>
q ��EگAD�l����"-��F�3w�k_4�5�M�|w�P�tN+=�)gc8����[%;�l�	pd���3Ow�. f����oi����1A�$�q��y��C��%�J�/�Bu�*�hH�]��	vt�Z>w�t��@��z�t�?o�0����ᣧ>��C����~� `}�8���O㢷$�A}B@��d@�Ͼlj�)`��<��|���<���sou?r�.�XC�5�v&�K��a_����=(��w7'��&A֔I�4?�rH�vw%�4�/���P�<j�H(�����QT9Z3���70%%3�6wqN��"ǫƱH�s��NDDբ�����W|�iI�>�L$>�gA;lh���x���>Q_W ٨�����{��t�`�Ud������B�� eb��7�]�l�)�bB�3��'���>)��u3ڇ�y�����h��y_ D)Q���A���cG���M��LH�j���MwE���8]\��C]�(^�Ɠk�#�F����9Q�"���!k~.�M�Q1������H���vY�z�������{�d�#PC>i�ZԻ�H��il._i�X��z�@x�.Ϋ�Y��5�϶^E&/>�N���4Ɯ�W�z�yS;@�� 4�O&ml�pW�Be�H~�\_R��%`�������5h:9�~��䅷i���3�roZ��p�pi�;�Q�'���+7��߸z+��7��(��;�2=�[Me$
�����<w�?Ɨ~l�@�<���pR��Iv��(�vQ���6]�o�	r��H�"w3���7�|_+!-�����u�9x��=��n!Tp�<�>�F!�����Z��M1���Q��\$$Ϛ⋲y��`kw�����]>(xM�X��`������:�E�;��-fy��?q\��S�	==���G݉�FV�~�{:�lj�� R��B�:ٷԈbeLН��y c����0D� 9��&8��Z2�@S�^jwH��N��pw]�[��~��v�����H����,��x������&��]�]��[>��q�(�lu�o�C��[c��)�{�>���w��A��80��ƅ��͌�c�W=��(��ɜdp���y�C� %#��]l�*�hXG������w9�;�9��y��M��m���*�*�̂'��h��aq����j�g��V�{11�0�	:d�A���Ȇ:�O(sN,��uYG��H��윧F�+٠;ͨ�Na�@�>��gh;��6:a��ʈm�Z0��E��ET����  N}5Y@*�d5Hk[��2bMe���<�eܝ��9��Z�`a o6	_��F��4�[ ��F��*SW-Ѱ����H�Z5jO�I���+�^������z�M�Н$V,�a9L�AEBb�g�Z��Dj��C�f�ki��#�x����"ȷ�&41{��YG��<��u<�ۇ��Q�S'9�r���6re��c��2�����q)���8��f�4W*վa�����V.���+��z{���n~9Tl%}V@j�F�����N�t������~7ܘXþ�Y4�{i��l�����B���I�`j��'f�V��1}��9���&����FO!�VO;��Y^��X��(e ��n��S1��ϺP��UdZ��a�Q��E!~C�5��(�&�5b6r��E�\���m�<�?�����*`��E��|%}�WYI�?�](cr�A%�V��@cV��_�f
D����	Af���H��ܬ����a�9�QzRG?�?���F��'O������/n�ǽFD��ѻ?���Œl�ыD�l*�{�f���d�3ʴƊ��\�ph
9�ٳbd��Q�TOA�CG�ڀM��P�B���1����ymO��/y�3>U�n��A��`�m���Fȣ��ʽz�{���	3E�r��ۚ~O��0�x[ :����&iij{X�2��Xj=E.�±+�' ε�%i+v���m��, ��`��T�őX>Ċ�\��<0D�a������l�����Ū�)xR
��먕�P�/~���{u8*����$�\!|�4�Ca?�;��@���n[�̱w$UwmO�������u,�pfj�w�4Q�WR���+~�t�(���7��tA�k�o������6���jЋ�#n���} ����N�����$X�$b��[@M���:�,���C��:�т���yd�ᘯK�n��͒��:��>y�=�o0��qc���7(je��Ob}�u��$6���P�co50�_m���D,(����A���	]����xHm�2$����v�R%�c��_��ɐ�߲2���''Y7��ב���.}�����*) Մ��䓞AE;!��:!iH��G�R��zo�A�s�7_v�c���Ȧ{���_�"A��C+c9Y����_�;������~�}��Qy��ظ��Fu�ک����a��H��J����S�a�p�D�%�4�d:�:�\	��b�P�L����ĳ�s��
&�M�������f:�qM��Gr�)L���/!(�J���y��-9Ǯ8;)�jS4��P�xk��n�*�݃�����:��oz����4z���]�t��u�O����3�|�Ø��nE�����l����F��v�8}s�4�C��BH|Ų%��wZy�xd�"�K��0��/��K�,Jg�C�Q�2���"���`s����g�Hw��e�4����%h������͝7�h���^g�C�m�������cX?�V�Ȁ��E�J�Ď�t��1��3qgSvV�`?��3��;G�<���a��X���@0f����y���1��}o54��A�y�a�!�x��ݯǐ�E	I������74�zz��"�)�������l�OY[H�W��*��6׮+'��VZ��Y����J|����l#v��ޙ���L$��"����+K]���D��q���_U!�B(�5����Bp�Z8�j�k.��+\�ܕ�C�'�e��98�"�b�XZ�����W)�2G���j��:o�~��_���!�x�DT�Q��K|ȳ�X�R��+�2��@���5`,�W�\��x�Z�J�8)�䦇gF��0,!���m�,�hpF��{$+*>���D{p�}���Q�C.WeЮ"��D�9, ��������৔�>3/��:��@+�x�R"�X�J���s|N�-�9[i���
n�v�>�R��/y�Q5�S-���P8�r��c��taX�S�WV��\�@�\��p
���"vT����!CN3���@�̐ӂQ�6Y�ӏ�~Fv)I���/+S���9�ʘ�b�f���)M	k�ҥ�aNF�Gč����ˎuy'�A� ?q�|��S��.��H� �N�:��N��1v�!�5�{�;��H���b沤���cS��|�S�˨�F��`��Z(����vԪ��g��3�TkgdPX[��Z�2��C/��n�˺l�)����*~�����ڳ���$�dӔ���ڷ:*����-�2�ȥ,�D��:�A<
'����6��ไK�Qxd�2r�j޻����1�l�O&���nq~$�-�V?�@&P�O����z����5�t�;��G��0�Bh�F�o��������~7�t�}���{��b�*%�z����`<2�p\ ��-�A7w����M��aQ��+؅VcI��иu�_�n�-F�M������)wE���pb晸]�2�
hNw:٥@_R��
�Rw0�M��L� �>5v{f����h���.�W���z��}@འ�9������h�[C��Gwak��%����cF4��8�P�C���®��At����'d&y�e���6%c��PM��1�O���3�M7ݰ��{5V*�����?^��w/��8�B-�;[S��������q[�o�}vV.<-l�wf�E�z���=��~?���@�ٺb��<_��� �;].����S-��H�'��4�����M�R�Qp���DYcZ�hhb�w�v3\`?G3Z�����wM��Hz�d��R���[Ǥ�s}�!�d52&�w�$�"���n5�|�\�
|ToNhЦ_Gp�I�[f����CʈR��L�ʖL$:�r˖�&0�!��z���N'~2۩ݟ�g��D���SQ2ܹ��{n��7�(X�_+ZX�;bY/M�l��	'��["�U�{Mk5�.JY�9?��l����V�QX�V����/��5����#��Iyruu;G�c��'��T����-���_Rߜ�fFs��d�ѻx(<��^ô��W��E�&�W~T��J�.?��KUU��������cQ�B)����0(��:t��ԷQ��:1R��q돛P��|���	8ʀ�)�� �ىA-"�9��Pe����Y�mZp�۟)����*"��V��G���"[w�Gg��?	���su/µ���+�Is���Rx�h.sׂ���9�h�䜘��~鰼�A-8D�O�[��n+�m�ޑGh��2?�Tz��Ӫ�FIէ�R��O���,��f��\�لb�Հ,��%�^��S/������㤿�ru��b�0=KpC"��������)��<�)���2uqLo���� `|�*��n;T��tρ�1���jD���q�z�>-�t2F�J31�=����u'�n��w���$�L�b
�4����>5Cf�Չk�BQ�$&�>�>���ݱO��:� 7����`z�f�h�P�DN+)�9�F5�-�4M�xU�3U����m�з�n�V�`�6!R�D�l�n�Z�`) �Ų����E��U.�	L0�h�D惈F��Ʈ�<����$�`��@�?u.5+y����m
W�.�D�����v 8��xA�=�ԙ9_Z9����p�=uu�@V���t�R�\!�~�e���m�ܾ�<ҭf֣e�9�a�[:m�5�ܝ��Y͊��#
6[�X�4!�*�T�_=��h��-�/����8����t׬�����=�~2-:��3�v�V��E���0�Q��8݀�"Pr�����HI�mb��'(L���O ���t�E�(���n"`�B��'+�M�x)Lf!o􎄙!=��E��l��[��Q��+Y<"'��>�v�M�{��@����\ՋhO������݂&9��5-Q@�D"�r=(̃�����1���L7Lћ WSf(�7�#9Fx���M�H��D��������S�@3cz��k�O��{5jX]h=)A{���x�������0�v�g�����g�_OJ�Î?�T�u�
�(<�J4N����QfЕc��ƽU��N��{�
�"��rɅq�� ��Ɖ� �}�˖���B]]���N����*j���U1�N^�'W�D$�yG�	S{9�M���<�Vn=d��e{��~�He	�"�X�w�t6��:*P�C��������ә8V���:gǨ*�!o�UY�؎q&c�+0�HVw�)N�		?����`���Á?�����֛2��Rh��� �L���6�}���Rس�U@��y�j�*�5��A��c|��ۦ0��KTs��%���2��Zd�MYA"<���P���2��7X@ʱ(�2�c����_���od	�k-��Lr�a��X�#���Wً:��o�K��tk�g����R����!�K��X��_�^�*��P+���O
h�K������[�����^<n�^;)�uO�b�*�Y%HBO�y+�t#��0B7+B:�y|��j}2�P�i�V/��8��=C(�$U����'>�����ft���Ļ-�3s�7�ԕ�����<eͣ�):�aXe��=���
������q�Di��L�j�$S�Yʝ��K������ 8NkH�`#��ym�X�!�v��٩ .�{�ΐ�%_�{1�w����t*7Or�G1�R�B��c�,P��V�9�Rڌ�f��2Õ��P�p���9#����N P�wk#0w��r*��(�Ŭ�O��Ȱ6�������)k���׺]�r�Y��T�/ʫ�pb4*%q�0tXC���{䮻��+~���Ω"�R���[�����"ɵƕY*��*T���I��7��ΓcA�iQM�]���@P�FOF�����
���U��B��Ě��eDH#����R^1@��;�E溴oZ����=�>��ǩ���Gz��!=;�w�������,�)�-`� \N�/Nv�����Uq�#��q2�V�}0�w�Z����d/v�+}+���MƩ?i�!z�J����ܾ�C��/D��?_zU�{|[�+�JE����@�Ք����.���Ϙ����Ѝ�3�45~���Ś��Mb�!_���a�5��܊�͊�2Co�8�[n� yo*�.ǻ=�h} 
�b�KD�E����ewB��g�#�e�d58��Y���3:p�E�O7���h���a6Dx�=p���xm������8���h.G��C�����o��?���-��y%ޕ����$t\Ͱ����bk��ݒ���#7X����?�0�5e>�.o�N�r���7D"��I��'�s�����U������h��k���|4@��r�f��J���1sMԝ��:]'ctPQ'	��ϭ��0�Q�4Ь����5<:�,��Y��Y;S���]�oe.�X�8����E�_�˅z��b�]߸��(� P�`��\��������@)�):��Y�ƢH��/��:M-���0zr�1����d��pESnK%���t`x'��y��|�^���
n���9�@&�J�W'�~�Ԅ~ĭ\
���r4,@���F�7����ʖA8��2����/N�i�ۛf�A-.CW�d�2@a���z:J:`�6���V�B��.6Ir�͢�p@,*`�g��ֵ��f�L�^V�q�Ri�lp	Q���
��yc�i��)�;���0�i6���4 9=т���g�>?;d�s�:�.�g�5Mj�E��0��]If��L�B�R���]�A�ȼC�0O�P��<�x�@K���'y<��J^��Zi��C��e����dE�3!+ �థ���NyÍF�Ț�sr�?�^��r?k���:|ak��Ű�'��.쀣�_�<�����c�uZ���S��C���iQ����w
� ��pF�4���=��ʼ,`�@ڒ��� Qg��(j;�7�R̲@���5�ߗq�,W
f<�����'z��� Q�*J�,I�}E@or��<?i,��4�(�q�w��G��������c��	d�X.�wԀvo��A��Nё�a���aW������ G�5�z�;'_��%�~�G�t!�,���-Ӛ��;�Z;�!c9�w|�@�P���
�E��@%,w%�mO���ui.,�J�1�:D��BV��e���Q�0�{����K�߱� �X�d��9������ iz�n �LP�q��*ډ �5C�QO��UaZ�ڸlj�}� �Ed��(��nu@V�����e���H�E�6	�N󧼜l ��]J�s�Z�\)�mF�/���7�T������Х�5$(��.\L�C�@���VB8Z�]yh7�_��-�t?�QK"�<#���?S�3�¾P<�Vu�#f�M�/��׌�W"�5:�-I���Q�vဳbY��M�c�@\�	$+Z�mj�:�q���T%H��w����`�ѕҘJ�J����n�24�㰃ьS�m��ʂ=����CF��9_H�l����D��`�25�s�$�V>I�c�p��w�%e��jI)LR��eL��nd��dZ�q���m�1X��4*=a��I��OAJx=�:v�Zuv��LPx�U���ϒr�
9ekC���7n��َ#�iv�
��7 J6���\�ԣbx�Y�9P؅��<F7�ي-��3B7h�z��4E;j�۾�1s�F�A�"��'��Q��ubԶnP�]'u�-�d�Y���`��ո!��q,�i�]X�5����T�`m�nE�O.VP��V���I�-������<3��k���z�y���߁р�_��J�OGL0$��$���]?��0��f�܃�o�� ���g՞�0bt�.�		U�u6�q(ġĹwc��v�&�Űw.��7+�L6ٙ���/	>�"UZ ���J}�KԖ�V�}n��#Мh���6@Q��h�d"^9ƭ��@[n`��jJ����`�W�e�&^�7��=$.Tx/�Ywؓ�R�I�G�w*�VT�1b[ϙ�*u�L��ɜ�}M��_��ĸK@��)���η�3��@Q,�A�c��@���@4�'w��(�kE���&��YD�M&a��p��`;���-u�/y��ʹ�k!_�a��G����x�?=���7�~j~�"�z9���ō�K��v?����e���z M�L^a^�\�zf�:�"��������a�;��/n���ݪ�~�B��_y�=n_s	�k��_����A�N���Zl^�g�OT��v��c�!��PzVԄ����W����y��+�l�cO?�rk��i��]�k����Y4���H���I�Z`��w)�/O�i�/.]�:R
���HQO@'ˊ�����!KU�s�Ϭ�k���f�V����&-sOD���PcV��z���ds�J������޽7_j!�a�qP�9�%�}�ܷq��؞��G���1T�F�z6� �ǉ1�w'�0�q��To�[��E�M���@�@�Mi��n]2��L��qf��)�m>�9e⛑߂~ ����FFx�:.q���K�������`>�$��Yz���t����ۘ��*��a����`ṓ�d�����b���lN@c�:Or5:�!�(�(��a��~�c���$��f���f�,���UC�[�S��0Vt�Cb��</�D^��Q�ٖ�B���ϊK�+T���s��7��q�Y���:��(�.��X����&?�oU���kJYW�NH{���w��3�6ZE �|�	_o}:�F�#M�4���(�͡v��x���%�׊���(���r��y1�SV���=[�x��E}�|�1�[��%r���L�c�%Ho�a��m�;+b��װMfPl��~W�z�yv)ڇ�qļ�R��a�'{º������"DB(h+�����8�Ƙ�c�3� ��e]��cu�$��.ya9&̢�������]�q6�9Et8(m��K�S��c�,0.,�n�W����2`ʉ�} �Hhd��Z�sh�,7�I���q�J}3մ���`���kl!"�t��hxy�����q��*����i�F���l�D�-U� �gbOԘ�Ȫ���N�p2��1���k֜/��f�gK�<&!VEq+b9W�}��]���-իJ�ܖ��@Ze_aɀ�@X�}+�pW���6E��k�5��4��f8�^�!��v�@�/$��KP1?|f��GPP]�"^� �C�Y
xW�*�y�|8�'|�9�J����f��h5�ߝ`dϬ�r��	��;�F?�e��g���aJ^��>�3b?~�rW-�%�L9J��љ[�Xtq�-�/Mdv= � A�҅�0�M��݇!^_�u2m��G��RR@H���ʔ���O.$߂e��R���k>�!g�I�UV\�P��lg�8>�qb�4���֮O&��W�ҪmG?��x&�?P������>�E�%��I��vs�n{��qo?xi�{��p��Y�^(2��1зj��fd^�:��{3w��T�̂����Z��DU����v_�o��N�<G��d4�zd�4H�ڬ%��3�������Հ /ֵ�y�G��ZT"�6gQ�0����N��?`���J��Rk�_4��O�O�����x�M�$�dE@q���ɮ�M��A�7>�����]��a�P��	-!x37I�9σ4BX����)k�l��� ׹H�O�Ƿ��M��u��S�,L�ٙ@?��D�Eld�u�%r�f18���5�d�����K�B.�*��Z�G"a���aA����.��|h)�Wg��*��Kt�;�d3,����	j}p�j�n�ӫ���R`m�^�/��afUσ|t+Ŗ�� �4��*�7���A����SBt���4�J�H�L��������>��4h}�`���;#*4���^͌��!���f�0�՘\1��j�������ۺ�}�\Bƹ1&"R�}g:D�%H��U�;��7�GS]a����N\i$�4����Z�|�n�s���ѭ%h5�#4Y���]D�;�c����+\��0�����BW�0���.Z������(lA.��i]��v�
�M�-��^��Gt�9S"�Uh�&X,��l�ϡ�y����;e%/���-zB�،p�oO��0D�3�5 wl�)�0�@7�����vyT,���A��٢ә�����JN�I~����%�x	1���D���:,�mA�ul��o��jc@]�����?�C��K�a-_�����DV��d�lh���t췢nc����O5�H���`诼?I�����(y�������l��oJՙ�٪����4��!t🮤}��4&)+L�,�V2Ϩ��Q�194Pi�6��!&ͥ���K6��}r�K	�cwn-�BH#82�ɶ�fy�<m�89�jB�_X
����9Lb|�D<�AÀ�Tw�R�8 ��@� I���0^��Ѥ�`f��jy����f"w���z1:uh��ZOcZrn8�8J��@�Y��8�P`�]Db�Fw�td��}" )�53>�%>�P�'����*�`.'�	�̋o�hQ'E��7����ڣ�<��n�;�ʐ-H �{՚����I����?�qz�ș�o:���oC�w沭�u���=��~��R��<_"��C���O���Yp[G�*�F�~<���@�T�^I�'I�^�X�P��&5��^�m�l���p1]��-�����ם*�/DDr�p����R!y�aq}��r;!*40��vfڞ�����Lw�Ew~��&6^��MxӕSİ߀t��n���]ML'���Z�e�
ѵ�%���b�����?kvp����q�5�-�8�N�Z��
�}S2�0����.D��n�ڭb�3ց����+��S���)a�bL�N��^ ���#a�1E���ge�U�6ڶﮜ� 9@M��T�y76���h��ᓠ衿?�Ȉq���a۔�x�e�����؇nE�z�9?�{j��M�f䲝�1��m��_�����	ӏ�y�͌]��}zԕ�rF>=�6ZUe�s<�e���Ky�ʎ]��&"�l������aT��7����{M�aT=�)��4�}"�;�L@m�@>ͩjO�G�͓��&5v��S�[�q��D��O-��IX��T�\Ю�D;(���g�6�5��d�:Y��=����Y�Ӯf�R�/R�&R㷺�5�.�<Y�ZU	X��>�ҀV�-|�����o�V���������9	:�*��ʲ�L�;�$����[��sP�'��
a�!	\p}��'G���3*��au�W�Ұ5��I�q,�+>/[Bh_mf����	�'�>�+��H����8{̎�4W��������j*uo35��g-d}�FnC��hm�� ���筱��.�!27�F���>,;��I����ј�$���T �XMP�����2��^4�i��Uh+�)�̹��Ha%�MU1�^�P	bb�B�G��m%�C�5�)���������	�XH�(�;�9�ęa��^Si[��P��x,����D��%`�[3��P*̞�*�|��8d#M��[#�F��&�$���
edŌ��<�?~�}a�$h�h�9�O�#�j5+[N����t>b��|�e�6��$�-�d���iÑ�X����]�`���#`S}�/�jsݯ��Ll{����VCNݲ�����0����Kd�_�I��AP�j�Ҿdxq��VΆ�9m��-C���p����a)*�Jb�)G�3���C�*뽥i�����/��f��x�1$"�X�/<u[:�Hh)+v��.�U��6b�t�%�S{uDڦy���*�|ǒ�|��m�� v�������x������*����Vo�	i<�� s��+���=~K�w�#��ô�A�z�n��	�[���0�����&�y����0����� g�m�f���y�H����/k��`�а��Ev��E��0慘ȫկ���,z�,V��G��u�[P�2z��0����s?�/]n��F Z��P�]��9!ߑ��D�Z~V�}�z(A�c*�<$��h29[N��)�~^v����}b���P��b!�֕�mQv�HOρ�
��Cl�ka���n������ξ�v+¤�%��-8�����{��{�jlV�H �_}�:�o��5.���������h4�T�B+����E��Z����|G8#p�\�ɣ�"N�Sc��`�ݺ�M�OBx�U�\Hm�I뻑�����Ґd%��V'��3��_��g��ԓ��z�صxS��B�b=9�W��D-�m�"e.�<�,�q?FI</��qx��|ϑ�w+N�ɘ#G�@j|""*��Uf&����R/[>�~ ��߽�����]�"��Z���YW�՞sc�Et�Aug��{�w��M��GGK�r3ÎV��{ֳ���j��H+Qa�������^k����ņ$��wN��:��+�c���`�s�T�(/��w �Nu����#|��j�-X[c���+?�� �!�7t;t@�7%DB���bdrw�Fs�<nf�S[�3��i'���ӖML��tَL���T��1S����xWcK�<S����P�r�A��i3�m�1��L1̍�v�[�C��%I�5��=�!��i|����k{&�TP��W'p��{"��.q>Je
w�dS��R,&dj�,J��j�Z��hAs�O��U�0�w��0mG�i���u@P�f��o�]�V�_��O+�O�&u��4�$�1�S���Ř�|���>�Fӕ@�V�E�)o���Y�]K�TY2h�	��{5�=��H��[IM��:�K�^}\6x��?/r��s�P�c�f�?�����>���ܓ#W�6�2�����St�>�x�~�J�dr��O8��>�W�^$�LWx4,u�(���z�2+�se������)%��F��[���H[ߏW��}_Z�:��3����&=�	,�.�W��i�<u�m�� ����I�3m^O��t]i�R
�u�� fZ���d��gjy�O6f'}y����K<>��?y
B�0]l�l0*n�Y��E����_ g��]$���80�B�z|�gc^�]l�7�*�.s0�Q�z8(����[���K��<$C��A�	�E׌K��rS���}Vɘ�*X���uk����/:��O����йܩV���_��30:�����=�U[��_�16e+\��2�%�3A ߱Ĳ��i�!n�R�"�j��h�i/"�񃫌e7�9Ò�̺���XF�D�z�h�de��Z���_C���P~F#~M�t�͠����`�����~��i.� ��p�O��D�~�G��k�M��Y�Ǟݑ��Q���h6���-s!^�^��"��fHԵ��I�u=��c5K��Fh����.~W�c[*MK��ȃ�����)�fA��6yw�m�/D\C�� X�Ic��9v#���!7T�M��)�+ �+EE9��*,�*w�Ch��pT�:m��1��5j�u]��=����0�Y�yK����4�֎���������t	��IƍA�Tmg�B���g0�'�l�e�m�p��l.'#�"�~RD�ڙI���j�Yʵ*g����(����p���7+�Ǖ�9�&8���. L��nV�g�E.�c[`��l�Tv�%(K�=	H@��R��$N�8,QQ[��JpaA@Kiz7_�>��F�
kg�5J՗O`7�p��Ó��ײ�)�Z	R���c�k�=�%�Ѷ/K.%֗�σ.�������ҙ�b���p^k��`�up۰�hD>W����w6[��5���D)��w�%���d�wY����Z2	qiT��u���pI�XG��	�?����pk��e����8�o�`����/"�Ή*^j%n�WcO�����a^Z4��k�_3̽P�Z Rb�T4�0�|�dDq���-Ό�j���50���'�K/����[}p�{�4��^�	�Y�q}�B(a��߶��v��!>;��U���t(f~!%5H��:�.A㑦P�ᄎD =�������/�}�K�B?�m���@]'V���Jٽ�¬�s�Fߥ:�(}	FRk=%�`��&;I� O�=���H����q�X��;�R0,v��^�ݩ�����pK�e����>\T7l�J,͚0@\�Bc!c����"�9$G���[��4��X�D���rG�P�yfG�r��݅ j��X�hĩ˞��
��lN��U;+����p��T�V������w��i��/ꤓ�T��[#ߙ�a��~D�pc�=�nٺ�E9�YdƕƵ�`aS(�_)*N�OV���V�Cg�`���ɇ����'s�ȷ��iE^�q��b2�\�f���X��Z��2��Ĥ7�IC���U��[Ǚ{�*cc����dq>j'�C���ax�,lϽE�xI	��Z�3����"^�LQ������/��&.��w2�_Q߉' .sp��3�T�r����EC�\ʒ$�Q�L���5�Ɩ�\B�0�g��@�2�K��ˢ�ü������!���w_�<����ʛr������	w��[5�R�m߾6~�݉EE&�,���\Ec��@?����n{��� �� �C�=���k��V��U�E2�(�����0~�Ԋ^e���?�-y0S'��l�w���JF�V����]�6|CҖ�]A=6��a�h���n�9����v�u�-˝�K��_�h~�mD��j��kʙ�6�t�X��!��6��h��(�%�"iAj^�q�-6b^�$��DdN��
`��.�GBm>Sz���p<��	��*؈�e�%~{�v������}���J|0� ;(d�-����3��tV"��;w�O�k�3}Rf��OQ;=� ���4��&�1�@>(��~����Sp?$��x*ϔi�K������XhHi��ɵ<?+�S3ǆ�ҵ︛E�)��>�NT�/�/w��^Ά��:g��0ѱ�[��>�6H2J��|��h�f��9�[}<�QB4ދj��F�c������<�6��[d]�X�n�b��Z4/���P����>�Ѿ�C8Y*��\��P�� �~mϪPu�x�4�����!?Y�z�
j��{]�5�1�b6��DF}eN˩{�
���Tz$��k�Qa�1*� q�[��4�=z����PÖ �D���/�+]c���rl@ݙ9��⧥�#\l.޷��"XQB� R
��i(��M��G3S�q���@G$2��[����yA̒���u�On��<�4W%#���i�s��Pһ��e��XJ���%*���u6�.�`E�=�qC�\>��X���B�E~}�OA �UQ%-
��ġ�t}4|2f9���\bv_W�d�mކ�4����,k����Q�l�k���-�T)�̕�y�U�dJH��g�5�.� ��"`>��#
���v쭱<"!}.%��[Wq���;Cd��mb���)�� ��H�<�9��ަrI��~Y鉶L��h�S�0*�֌ҡF4���݆QD=|x��ĺ�gM��"��D��*U��l�{��(�z_���օI�L��測�glz�k��qA�VP3�$X�(E��y�����g7�䥽X��Y��Uh�B)�H:|JWRZ`�s:IG��*��Ʃ����mA�/�d�o(�'�}и�k7�X���4h�tD-��1� l�Wp�y|-]�Y#,T�����Z�LH���s���s�����ꊍ�3��xr�|I��ȊW��E�J�����2W����������D�P�jV鑫Ջ�)��J<�i<����9Y¸�l[���e���[a�.ƨN������>�/e��)r|�Q{(�AK�l��sNt����ع���=����g���]���S�[쁒uB��	������%#R!l�s�>�pˢ�m�2�[1��-F��7s���w����Ub��LɈ���a�3�ЕZ�r�`i�W;tB3��6^�`�w�c鯀cf ��Wi��݋>6B�5�/��4I��*��M�rwYgak<���Z����ʛ��}�)\́1
�ǞA�KaJ��7+��l��H=���[�ȃ���W>�S�og��Tm�z$�wiڕ�/�cIY��@iЂwS����L�ܙ�F����
��$��S�#{8��|xDb!]��V,a֦��#��%����5ؙ�	ڷ�{��#�J/�65Q�0~�b�ן8r���+��m�ʭ��|�d;�-���R����&E=M�	����Pڦ����+�it9),agJ$��lS���@z�"-�f��2R�n����Y9�8د�jOw�W�SO��,�)��#�U)b��%�s2��e7��یY�^�b F����08�ޓ5��
؋7/��\C�� gt5�y�g~R���=nQ$�P�ۙ��'�\���W~ג)��c?h�WTf�*���G�q�A�<,F�H(�X��ט��bm�b*�f��U&m��r�Sq��T]
�$Ţ�p�c?��)ڀu��Ev: ��Վ|H���}�뫨}}zm�Q�4kx�hGR�%�y�0ӆ�w��7���K\0���cil�z9S�me"���!�1D}�� �����oP� �I�db2o�p��Ѿe���x�nF	�"�&p�le��y���x�ۍ[w_7r5v8@�(U��a�ȡ���XC׵ S)w�]��
l��@��0 �O[sͿ>��������E�L6ƒ���H�Qu��f}��|���(V��l�-�M��B���An�b��Z�y��4ݦ�)�Ν]���͠�����|�zX����y(ԷI�y���~{#���-�{�F�(�d�}� "֧��Qpb��~��li�إ��$)m0�";	}�*+��2��sS߾�g�a|� 3�l��B��@C�Mx�J���|�f!%��mMgW��\kZ�Y1���F�~��i�����3������ȘB���TR<o?t�$a���}��5Y�*�[ h��?�<���׏C�=5�/k�VB���S�-����v'������&)���q��cA{*Vm�mꚆ��;�-2�"��z��_U��1��Q�\IA���Ͱ
�,Ê=�P�O�=�&m�5{Is	|��g�bfI�ebKy����d�����Z�4A�K�H䞄�- 7����'A���3��[&I~l%��Gl7��+�,ۥJI�C���g�"|̗�&���~[���6X`���l]%�Χ����j����\���l��+.t��d�rF	MN�;�]�碃>1mv-�M�M{�>6b�Ʒ�-�)i$�6��"�7�i�e�n�C�o6H+����t�7�LE��f+��Y�@��E����+��3�nj�0ۦ�g�s[����n��p�~x��<�[�C^\�u�w`�e��~8���*�_MlZ�w��Q���V�w�,v��r&&�4'�l@�l =�\�y�,Q|( ����<3���O��p!���63R �OmD9��6�Oi�$�r=��"i�8�u��ܹ�zi_��T��j6ҩ�� �#�K�\����̻H=&���(��U@��;��(ճf)!�l�a$�$��Z�\K
��Ti-����G����Y&�	N�o�uS��Մ��)HS+$+l%� J����H��5�����7q2���H��>l h�j������E��E;���`�2�k#ɏ@�zlLL� 7���H�:����:a�\j���hՉ��g��\	ǟz�y)�]|�UU�f���o��C���W��)�)���r%�.�Ҁ�+��D��p7�ۋ�Uz�t<ټP���Oղ۹G��9�'=s��4(2��+�3��U�yy?s	yG��3���(��&e���cG�y��A��N�LMI�i�J%5U��zr�<��4t����E�0���u��}��gD��AѦ�7N�,�ŉ�jA<�d�����&' �gG�2�4zQP��U��Aa�u��ܑ�=C�t�� mcgu^�����a.�Jd�����k9�S�y��LF�,���Ƀu�,}�Ǖ�Ku
3�ت(~����	H���1%��}ߨ�n�9����|O<�(f��L�u����=�* ͇�q[�����Ke�P��'!÷ձ�'5�K��O2v� |k�]G���]q����C,����˃ږ�i��%G�C���6���]�[J�ӝ,�A�J�8���k9���&&��]�!W�%�?0��Qc\\����*�2U��6�*y(ȹSԺl�!y�Ѷ+�<��4��H����!��r��$�	d}`�)�$�����v��|�$�;�_J����ș���1�	�h'��]:��b�������G�W�k��%��I�e��G}�%W+��!p�p܍�*(l�.�����R�)�_~���`Ӥ�{��H]!��[T���ҏ��1||I�9���/0�Bj6r!�P#v�6��hy6�@�ak
���/��.�ti������A�g�7����r���݈&<(�������*ȕ�2������g�}�g��0=XX�0u^�!��?��M��5_���ɪ��1�`�{�b�M�KPs߰�����q5?e��\�S>�^Y1t;8z+<��႑F��D�}s�ߚ@�^���KR/{��n��ن�V+�Ҙ'�L-f���K�a�B�|(�Û˧���bW��>��S	�4�E���OB�$�`4rL���2�����]4�ݻ>r�S�3�~��Έ@<��5.Gj��{���#��pRN^[��3� y,p1F�!?p{��?��GO�aL���&��b}��Z�U���5���&8+ZG+�������0���Z����E�{�6�hn�9$L??.�s�SM����
S��-A�����ݎ�$�����u{������dMhgz��2�<P%�i^�xRSդ��\�g���Ä,VUŊXЀv��ׂϰog�]�6#Z�<��Kd��N�b}�J�6�2O��t04I�e8[��Z"�x�E�Ҳx�@�gQ�炙�5rcD��^�.����H�C8�A(T�|�ߩkm��
�V��EL�I�H��K�C����T(_K����1���a�)�Y�==ܓ��d�Ć�E���@0�{���Mu�S^(�C�cF�*�"ؾV����=~E{m�¿������T ��b�@�Katf7�3��?���������o��ݮ�2"�.��6�����=`Jޓ�Ae�
�D��I�-$]��K�!w��~M��}5�gF�r�����8ٸT���N͠ʋ/?�*ꗢ�r�;M9Z�o<s�m�7#o����<��un��`�d���ߺ�#�����r�������x�,=^�K�Jݜp�(9a�ݹn<*Kz�K&A���[t,g���@<?v�bؔ���nL�Q�gA��K�n2�z&�g�'�z��%��~db�̈��\�B8C����k(`keg`�T��
>�o��k����/�U�(.�@��@҈w�P���p��.](��N�� �E c�LW� �hLx�sc�h>M��ޖc�#�2b΁m4'�Fg`o���v�(�l�NX�Y�*���p�4@sC҆��j������lf�8@p!�)�������{����Z�W��@��X^�(����X�s\��g�E� Ǥ��UZ�*�*��oi���ʬT0�Ra�:��#���w���a�Mԡ��~ܝ9:���m!�3 FNq�D}�1��_rA��	��+�a0Wh-h�rSwW���y���3��T�G�S�v»$z7�Gc�3�N�!��G�b����M����?�j�;c����!�|nB\�euΎ��U��7�9��ѥ{8t״aL�[��C���Dsd�Ί�LcE{�<)hΣ@Xiy����!(�tV6��y��`�*��f����cl����1AD�ȶDC����;��(���5T�2M�2�b��2{N�{ʍ�ΥA1�Y��c�!=mP��R�p$�a����+w�����s���� w	x�3+PGӫ��F��~(���)�F��ǲ�}j
.�h�~d��bu�~�(&�ik�ʹ��[�9����0�(|}��ԇ�-��y���kEU�aGG-c�Y^���g�����#������N��^����������nf�Ź�f��Gˮm��Bhk�Z'Ώ��w#��g�(PU&dnU^7m�T�+�>;��|ǘ��膈�/��|�T^��j���m-�C~���{�6j�/��n.Y���R1�ơ����%�ʬ�����sӀ��9QFx?1Ҁx
���7+��`Zf�s� ���_�_�h
j�c\�@}��mI�\��PYР_[����E��B9C1����s^h�Hl�Ȱ�DR:2t��7k~��ݴ2MQ���֧z�+�}a��
'U5��|q�4'O\@X<�����z��F��
�p�oX��5����K��.i����So�m19w�OP� b��I+Ō;��R�p˖���\��������$9���!��ʀ�O�4�ُ$2㚁���M�]�;c�W��r���4�<�SWR;������:J'�0Q$_��-R7a`�MR&��38��C�>j0�]f�6,?�j<� �T0�J8��'&9�1�oN���1оM@��=]�fϜ+=vu���6�ԛ�[U�vζlYc�r�5D"ű�_XKg�}l{��,|��+��q��\^ݶ�q�O�Ab�J�.��t����F�Rr��y��1� �V��& }��No��6�ls��C�>O*�A�?�}I_��������ZG<3=m�G���a��?Q�0����ĳ�A�]`�IPZ�7�|�p<��_z�t㾩�F���������^[�#{~���|
��TP(/�KFU �&0�����R��b�v1uqx-"���fD߮����^�tR�z$�K��|��١`�n}�?�L��l$�� a�����d/����0�	Dz�P1�ǆ4ىЉ`���{fE�}ѭ��,R�ڲ=��F��Ю�r	6���ɠ�� q�W�]뼫�a>23�3�|�sa�:Z%f�toqC�ߡ��/6��t��:�NOj�Ǚ�aڶ���i����eS�D�a8�ef{#>�[��0Xk�"��Hc��� Q�!�������٥�h�G��W����ҥ�O ��#�QJ`$Э�l�3�%#�G~���Q�.O���l�~��`�^p�0�����Ɯz�Ō �H.��IPx��M�ڕ5�%����o�g���Қ�V��S_����TBs�[�Y�.���F���{������P�T�-�dm�|�(q��pRI�.6�;��ro�Y���av���+	�|F+fז���0M2�����"�7Р�m��+z� r��0��%����e�q�fU�II�q6
��Z�4�8��t`���e�f�g��=�����Ը;j�I�K��a��D0o��(�� GKA}�&��&��w-����eF���p����w��B|����^%(Jr�!��A���Ob�K^����m{���}�2�9{J�jB���z*���YnUWbu��70H�ل8�lqyp/�k�Ϛw�r,�+	�	�X�^\|uM��lB�đ�A3��n�7-��d쯻�R�U3D����p��Ӫ����9�MO 5;͌���l�y�}1�|~�(-��XI$�y�έm���LU��Pae�?�y�s�sp��{�̾N�L����leg �G"���AW���'�{+i8�d1�q�i����꜅�_�cC��U�}B��">��u��#40xw���Je�b�i3�{c�2�`7��օ�J��~j��$�e��\aHr��)��
��C��
l`�� � �|�s�����G�ۘ��eW�W�w�>R�hr���!e��2<�ȻKy�y���}�w0(���~�=�|�Pӭ����\�:��'][��:x{p�t��~S���&1����n��y\h�u9�QO�	���#T7�w%��e"���H/
�Y*��^3V���6Lr1�+�e�d-Ph���u(�=(�f�sx%,�&��b�>(�WNH;��%{S׆���ޕXi�<b/X6F)�
_�b�m�`�CGP-�ݭ.DI�'��t����qw�\T/����9��k��,0��_���M
��Ḗ�d V<���3²ͱ���\>r���(�^D,������3��F̥��s��g��T>Sa�\�d�5w�6PG��5��#�DRG�귍�ʙBXV`�v>���ĵK��c� 8v����* J\�w=�ִ�<YԆA��A��a�2���fK�8h#1wH3���X�ߤ@�\@������C"~�����g�e��z �,��4�F��iC1�EMۆ{���E[l��4��m�5���y�7�:�����]3�6O�~�O�ݦ��E�&,�#��h��YM���]�޺тL����Tqw�5E+&�p)5�*1�d������&b�2j��t�P	����_���[}���0��+��}m�����L����źh#�g�n�e���X�
7z��o�B���W /K�2]�%9�+ՍjT������`#k��'�9�9�5P*��g�'Yl�����y�tLX&�v����^�
!P��rG��	x,b������.6�D6Ll�T�QW���M�_��'���`\��B׾�k,(�3�v�����e��ëc.C)3�rrR@�Z��{�7Ѿ����6����K mi��6I'�лj0�W�5Q�=�y��7��	_�)����Q�Z	QM����+~�+��O�m^��DN�޺cJ?��'4-<��W0lh�Cwv���ٱ���V�'�/�=�:p���)Ě{:em�c�OD����e��v�g$B��z��థ�BL��5B��4O�8���E���QXFFKF��N��|�̬"�mykw�bg)?���M�IMG����I8��|�Q��ˈr���I�� fDG�(bw��M�ӼE�vΰˏ���=)QAЕB�,���xX=���X�]!��� �8
0�1(O8_P埴Y�	��_v�.�,w��R�![�:X��K� �I˺T*�T�a8�aA���2�͂��#�(�|�R�k#,W�;HfZ�A���x�>l��=K�Q�8����pr�ۦ�[0q�w"n�ao�t'd���wCj�Ur�\��f�.S�7S�9)z���8��\���&W��Q�`�V����u8> �:,'l�"e 3��O0�=��e�Ӂ��D��!�L�#;jd1LW�3��c.���wC�܎�������7�}�&�?6�_̷��p�[{��yG�E����Ӈi�Dh�/:����˳��NL�K�i5M?e"��#wW���\=D{lJX�v7�h%�C�<0�"�d�����g�]������r���S;eš���Q)���V�kA�y�Mq���r
F[��]�� �Y���2�0
������SSG�f���A�Q�d4R<��$�9�!=�җ/ܕ�?�Bz񻒓���ņ�FZ�f{VjF�"�z�Rб=qz4�P�=�*�ɲX���#�*��Gd:�#�Ԡw�(�`�r/��Kk�xjS��h"��b��VG.K��>_)%]�ɠ̙����-ٚox�Ӟ6_��3n�8�_���5�綏�$��MI~N��3���1�jw�-�,}�0�Vp��ã�/u��gZHzzF96��~M�$���������P�#3=��\�����K�G�2�1�V�Bc7�ϼ���rɃ�5�K�l�g��� Rܤ�`˙X��BH��t�O��ս�&>��q�e��6�K0�"��e���.�Knw�;����_��J�@)3�+wܨ��U���hǪA(;�LU��Z�j�Vd��U�~�t4�U����>O�v����u�+ X��.t	V�o�58����*;�S%m���A�<�#��QӱX ��$�:Vs��f��8%(��L�:�@�͚�����s���V ��H��e� ���Ӹ{$68U�Ǘ�E0�L�\J6k�5U�(@�B�|��<�\d��:PPV���%����7����f.J^���ԙ��'�Ǖ�76�=�MFq��S#�.�G�3?�a�ڸZ
�t�9����yY�A�	�
el��@��r��\����}�3��1���jT�ۧ�?sU��Jܤ�j��v\��և���C)1S���@���e�ߥ�_B;����W��ܶ���1q�����?�떋p{S��������_������7W�oAb�}��ãj�8�XIL��Ώ��?�9)7�%O���w�:髽�w�[ɶO�<�F%8�JlM��j F����FP���q����%�s'[y�Ǖ(g��r�`Q�/�|�����+&2>�Bʝ˹2�$3�j�b*�B��d\\�����|��q5�s��ι�K�s&ʿ9��w�1�[8�S�*
�y�U�����'�a���'��$[&��V�V��f�ˣ�\ow� 8.�*DOy� 1�D�������((�!�x��tG��^�ޭ����_P��_��[��@��]�DU&	�m�[�*�)�q��sG�f*�Ǫ+����D�o��V�AB �6��![B�cμ�#��W!�7��}@/f"��,�NA���5��MB�3�R+'����/��Qx(��]ck`��{�[�$%x݌� ��\z[��������`NP'����4�u���:�*�z]�M~�Pjfə|(TσF=|ܔ��|����:�w����m�za�F�58�*�?����o{�NQ7c4�{���6go� x��h�xԔz�f1���n�45Z1B����zȂA�A���2�k�F�*��]�%���H���g+d�j�{j>S�&���S�<?N2�>Q�q @��jh5���\��6*��O��٪�F�}����rP˜j��D�o��]���ar�$┥]_jc��똃��������x(3@���"S1D8�T�ٖ	�4�{m�\#��\�ij���n�e�'�)���^ϵ1"��'�ì�cM����:�Ў#�g�4�ߵ�� [�ksSo���1WS�L��10�Gc�8�#h>9O����\G�����+�@:�*�G��g���"d '3[^��
������{���ۍ`ScazMw$�|1����g"�����Y6G6���_�
O�1 ��0����;�jM� �
i�G������و��bw{x����F��,Z��5Ҳ�[�E5�����M8�Ii�^�+���/녈⋍�y��@Qj<*��;��
s+W�Un��&���� ���������
c(ٔ�g�˒7�R��PyV�t��t�{%(�-_�ܚ5[�ls
��巌T���|Qa��r:���=��GR��#)*O;�z�A<�P /ᢐ��yi���(��!�VZl�j9���̅ՠr%��cA)��*�Rb����='A3�`����t��A����ˎ�gr�18<�����ٍ��(�?(���n�9r�|c���9�Oyn8�2s�0ZFd���`�i�muڀF�d��(�f	l��k�q6	�d,2�0�����.�ݮ`q������^�Ĳq8��*���q�w£�)P�s�ֲ����1��G�&��{��n,מ���M2�6���ˇUX��r���4���[ʴ7�z�����K��`��F�0�������� ��ދ�D�ОFf��C-�<go��_N���s����P��b�.خxDwJ,N�Vu�J|�C�ƣz��~���`B���0*��X�0�]���N�"7�qt���/�	U(���鲡�NfN�R�N�@�>G}m��+K�t�&��$��gh�630{j��/�6��[�)�լ��Ó���y����p
N��F�]:?�b�ے|q��mN뚉�X{�6(�v���� m�� O��;!���M(i�W�2U����ˁ�%�Z��'�1&y�N?����m�]��v^��puܻ���'1S|��?tO��Zv/��(��G��9Ӷ���/�S������=����eJV��\��)�)���J% h�e䥫q�?��mBV�����~;c�g��s��Gq�G�z�F �>�U?�s�0)�(� =Y¸��MS�H�{�xx���6��9K0���se��!��zp�m+���4��z�y	��}��݅��垐l��)����aU	�葨5_}�bZ��a�w���x)��W��+T
b�u��W.�K��M/�z���_��2`�s��'��Bl�)��V�J������l�TRZf�g{���l8�*��{}{�s�J�Rq�����]���L�wWPx�B�̧�h���>�'�-�8����0�nF2�י�aZ���L���PxR��c#y�I�_�6eCq���\��&�o��fq�ҥ�c��~��Pc��Ə֢'<������G��o��a�N~�_b�8��z�@}*�7�7�&3j2��^�B����+�	;t#����F���n��U9?Q�*�|��"-�ǡw{�@B�Z���$t��*EDS�f�3��zi���3���z���)�k�q���(ui0�W�P(T����uǣ��$/�-EA�P��%[�օ�W�0inF����
y�س�AITө	tPZd'�q�1 �"�lL�O�2q��O�5�9x=�gC ��T���!"�rBIt,F��Ԓ�oN��&x�7�����N����<�ѽ��N���R��AGI�CI��h78�_�h�I}Sj��}VuuS��"��P�$��`��9�v��Hd��|\�5:N��ꅂHo�;G��71DJ~X��(� ����|�-m�%�z&>��o+e�މ�T�drP���ex��\�q��/]�Q���I�w� �//�/pGC�o � �/����$���~D5B�}XT#���;銒�aH�d'��>l�s[�$a0�d�f�X3 Pr�d��w�)���V9��g��n<z��Y�~ޓ=P������ w篛���+s�{g����R�b��Sm?���\#H���'Ks�(ϳxl'Bg���楴["V��~�6b����j?,��c�����f���ݟ�!�~��z��"5��jk�(v�t:�e�k��- �.z@v� Y��y��C�����fµ�߾pR�d�R�F�p~�.>{�.W9��R�p�gw�-}��8��)���51�ЄT�d(gO{��L����Z���c��/ڐ�q`
��(�B��L̩�>���az���u@r5�]�:	TXR8��p"��a�޷��ƒ�M"y�LR������G���������������=��4C�
ذ@���/}'�$���ߪ�ΐ����}G����t)4"'a8>^fW��_���9(��f�0�a���}�y���X�z/R��T�S���Mж��������ـ� G��f�ԉ[����\gP^���|TC�u��rV�Na�EK�S�|���#�0��n4)5l@����-H�{�y|�*<�x-�ҹ	Y���+WK�7\)ū�C@����|�}�za�L�U�k�t?�TM*�(�M̌���	�cV��!��x*-F�g�qs_N#:�(�+5�A���t���$�p�u2�Y��?w�=Z�ՙ2��u�G�[�.��<Ѻ�/�s��q;X'�/���k�������ڗJ����6��ZG����	�,��Ɏ�x�y*g#Y5�Eq�H.T;b���-���e�Jb삏4@?���K�Z��7-\@�*�r{rĴ�=��"{�Ѡ�j++�P0@��v��=J�7���c���:!f�}�"�$~�D�H���0����V(�ĸ���"��Sӱ�u�c�˘0O������ၮ䋀��8��ޅ��C�3i;�9]��θ��1>u���6���sB�R������ϷD{��(�q_�����s�u"<oB��W>�-��V���$�L�<�7���M��_Hx;��4"z�U�cTRFF�������0�쑓��|�.��9uԵ�6G��z��~*���n�=o��΍����j��4;T��o�οRq���?t&b�~�:�����	��KKс�
�����eb�h�>�ǆ�3:�:O��Wsg�����
)}�&�m��7�)R�K���m�G�������o�ҩFf:v�?��D�n�5��u��6-++?횣�����A��\�qn,ɜݵ��u�Ƀ?F�2
?�:P�	�	�8J�Q��%�` � pp�g�2Œ]E
sebM-<>(�9A���o�a���O�&bj�=z���/M:l�������;n��Z��`F�W�3_�P`C���6C2�	� �s ~�C����?�14
?lE~"Y���9���z���p�a��2t?$���Y�yv����ȅKf���A�����2�SI�/�g�b��� ��+��M^�x�)�h��V�F|�$loCar��KK����t�B���!d��Q:.��:?���T�f�ƫO���R�z;F[�,���z���3L^�9� �qz}���%s��3E�mho�lݬp���0TSj���i�+�C�^���9C�?2T5�|�'���xǵ������QP+�ȭgnK�i��0����9%	�>TD��[����"���,�������/ĞmB��%g�9�\��K����^�pm�X�i
�e'���K�Le|��C{ep��k8!��B���x��]��@-!
_"�_g9�������<ɟ���6���B�����(JA6̅*�5��	��SND�)�N����v���(�e6z���Ae�K�`#bo�!���L@�O�J!����Aq���&6���y����Ԅg7#O8_�UH��T���)����(HbϽTO07)��Ɗ;�蘬�t�ൟ\�yY���$��xs�����ph�D�k�n7��LX�sC����b�P��@.Է��\X�J
���U��0}qӅ��	x�x��!��n�N�L�t�Q�>�c��q��>2�������;d/Cn�N�킜>D\q�,'����\OW��	/\��t<{�
�����mY4�=G�%u\�-���3DhS�9�[���h*���Ya�oK�6���J�9p�p��A�٢�4������$��[�R`��7s���]�/u^���%6�r���CrT�>��]4�����!�%n������r~�5% ��x�5�D�c�{��mEi�鍾 ������k�[���"�+xǒ��^)����qM�K"-o�Qmdφ���x�i���S͓TD�]�����J����%���{i�9�>)����1��3ù�zT���@�8V�S��U��"�E�9C�\h�/$7�־����Z5!^��Rgl( �����I�m�-4�6�1���6 ���&�_�]�+��s+��	�vH��(�D��ʰ�r�jvu���IO�ރ1;��9tN׫^Y�MdZYpE��/�J,{U��^:vKM?�:䛘�e��`���H��OR���y��q��\F�)_�����f�I�F7���*TU�=Ф��hbQ�*�3���S�x�˝�TAǘq:�dj�D<�TNG�Nd�����b�8Ky�JljͽE\�xe��(G�r���a����Y��HJ�y���e�ۋP���I�@C�Ҽn��; �)�h�Ã��r���htT�(�c���^rTRԝʫ	�[<�;�?�f�k\�AVFdH��sƍ���؎aX���]�024|@V�! zѯB�\�E+Oj}��1�����)-sG���\�v=���WV;IH>�
�r59���0�<�c%���9`�|�������86�*��{\�ٕs;�^`�x������-�׳�se�[b��5��Ob��I�=��6���2b!�!\3���<�8��2P`\�nIy�m��rB�:a]�J{Ao�Je9i��n-Ij��6$�{�w�I��$ݒ���c�c��0)�L������+��9� ��Qw�&i�o����>Y.��V�t*̩��v�0�:X�r�eV�:Q��o��_=gC�䥁�>$��k��7"\S��ƌ3�Y���N�sN3��#�|�a�#[��TA	i��_�{|���	ęт�Yڅ�ED�K��y��ϽIry+Q��ӻ��.��!����I~('����� m%}�j���'���_���0Ջt��4�a"�z���&�E���[i43�7����w{�6OKzR��m��G&�
 J#"�a�_
�>ߗ���?
L���gC9M�wՄĸ�C.͍�s�� 3�m�`���Ǘ�h���XHUqP�]��/�\Kp���] UQ�,<`yAf�W<�6qiqnr!b�r��cw�s�*�^�F�!���~�:?J�) <8�Nԅ�M[a��"0>"�%硠h��u\� G�C*ೌYh.�T���L��� ����{�11{┬��Nw��e����O�Ml͔3WS�֔�1��q��`������}�uG:ƌĪ�|��u��O�w�[%�5����������
Ԃ���Y ��'�(+V[��4p�q=_��U��,L��2�E��#�/GNˑm.{d<�1�}�P���d��p'�Mӟ)�������ک���0���� ��`fq��4� mD��"���MA�l�J-�*[��W�)^����J�g��tkZ�*7��QkÉ:㎝q��?��V�l��U���̋�䇁�}�
���b��rvo��U�$��Hu7��x+An�L6�'�.�UU뉦��Jdt[*Д�!$$��;�mͥ�<�����ڿ�sw��|@�[��W��k?�T6v�t��&�
�Uv�����`5W�,d>y�ȕ�G�z��H�=j��F	��������f|����N� (�)���G8ó�9�k�8�_��~�e76�3���a��Z`WF�7�sқơ`l�z����A���;�ae�\��kr?���8��u?($�|��Q�ħ�=����N�����c?c����>3�C������ݵ��2����s���IA 3,��_�0Z)� &�	�M���"!kyjY
���G�"��V=�UA���Fꡞ����yؔ�"���^�N
�Upڈ�[�{����p������,��xϢ�7�P�N:Sn�ױk�(���X���pD��K��5L���ן�}�ٜ즴�s-o��qJ�5��#�aH˨����\ҷ�����ފ���Z�^N�0u����ׇݘ}�F<ĉ_��c%�Ɯv��}2�<�ev�S�y�~��b�lIhb�-I���i%��`�����
�lz���!:�t��
��5��a.�6��_�$��t}�m�!a\�je�Q\k�T����)t `O��f����d���d�� A���f��6��~_C���Q�("\�p�$"�?F��?W�7,2��'B�suMn$�m�Gq��+�ڤMC����yɯ�V�	��j�M�E�(�"���W;3~� W�`T��'�	IS����R �U,�q_*'"Ê�F��,���5�ul�翜�}�G�= �o��i����Bf�n�����6�p2P�r��s\{:�v��!�K3��ٟ��$��At�$e��`r�C���[����.a��B;�Xd�Hl`��	�]ݝn���Fꮭ�<�����)3\��v���}�,��>)?D~�P�t�����<�P�mt%�A�p6D!j|��PN{0"��5�쭂V;�����(IN�f]{g�4���B�3iI*���ڦ٩kx0T�Ms�@	�u+�)��n}���м,�O�O�xRN��FX�Z�W�r�h���gz��n�j��m��:]Ol�d
H�p�.1w[Wxd������7-e�a�i����7<r�+�|�D�H�u�*�챦��-�h���/���Z�¶���aؘ�M]k)bS�gԻ�Ǿ/�M�z;S�nO��Ӥs5�����]�X���BPc	�̀���C��&�Fq�[i�:R�B�&ÊȶA���1d�}�0�ʕo$�՗9w�dY����:�T��8����vo����J}�j[R��sK3w�TV��/P=���{A�@��Zx�	J�o-jj5��Iq%l���d���n�|��x�}zf(O���糯%n;��_4)��̑��E��0�r��+�0�KϘֲB�N�V��̝�a�u߅����y�I��=̧��[�������o,ݝJ|
\��K5Z�h�Ñ���؁�Ҩ�/|��!r�^|3v6q������sűӳ���wEŘ1���]������a��8@M�oۃ�;K��c�M1��e�򘳩p�Ќ���.Y�۶yr�D�3cdJ�N�H�P%�h� ���~B���Ej���Qe9A
�wiʆY�s�0sVZo���nr������1��k���s}&+�q�W��#�1I����������VY��+�v�q_�inC���^D�+��o� ���i�Hsl1�<�Y&�*��� ��e��F)��&-���q��v��dڽ����B��,3�^�k��lWJ�R0T@`f��t�fbpw��!���(&D�&���\���w��f�?�-�*.m�߇+�O�h!�7v���Ǿ��n�`F������g��x���?[ԟK�L(|A��,�(��,m���$�Lsf<��V����L�T��+h�S�'k$c�3�Q���%�8#�� yQ��9���+0!�d=wAv"�����~��*�uT����iI�}�Y�C��2��1Ơ�m9�����bÀ��y�U:�'@>@ESt�&�q!�Guq{h\iD����,�D ��l\H��h�O�	�� %&���v˨sO:�䊇h��%x�&9�	݂�I_�Kݤe3w�u�O����&ϙl�##t��!v
�}�*�=�h_a�q$�Dԗ�v�<�� ����0�pn���Ls�K��G�/�Xp���sғzb����,��1^�4.��9��I�n+�LjeHq����`LM�Ӂ�/� $P_F���f�Xeb���H+\Γ��A����tc%+2M��Ɇ��GCv~q�c�/^n�V��a�.����E0���/wy(*�� h��`)X�!�C�q)X�+��0p����B�VGti��q��S�-|����]:�܃����t����Q�^��@l�CX�-��sDHM~jw���%f1&��bu�����޷N�ob���U�L�����g�j}�k�V^�b��^��˩�I�Z|���ؓC�K	m��w0�H�ĕ<�F�I%[87�~(�F C���l�y��
��nP~=}t�s:�![�PQׅߏ1��$�@ ַʘoLcI���Q.��hv�'/�L�h.�yX�~��mR@I�A�ꇍ�,}1��^)�F���s�`7���}��� 	��\iv(�wf��bG@FCy�5��v�g����о�e�
%��Q���K�?H�pRy8�"vrp�<�����V�"2�1&��"������>���P�`�b̦C>?�pCT�b��֎��i�F�=�A�W��~��r���sA�S���q8T�ט�T��xH+tL�SmZ8Ӳ#���A�w{x�ZSZ�ߪ̏UhZt�U-�1�N���3��{�]����#iU��+����Č�9�}Yh�i���l��\�a0���7` |n���qtB^Qvj��Ҋ3bv�l��$&�on����gqK$�\�[�}�(*<'\�t����s=_:ԩ�M��v\X�@��!�7�-��ɾ���vP�N-��V݃��*}ѣ�Hj՜���6p�Px~Q����	O��&��HA0p��r�Z�S-�Tv����,i�Ea%͛�����E����}�ѽwW����IbOA���n���Y����f���,��~`|P�07�Da}�ZY�j�>.ܜ%x�Lt�xU��&��)����Π̠��t � e�a@>��J�����?"�!�˳ЫJ��ⴲ���C_��2�l���]{�E������,}�"ȇS���g�ʝ�X'��W�퀙� ��$�h/�J[�2��?��V��Ul�ӚYp9bܻ}OyI�ݐ���tv��#�h3�({q�7��}�O�cY��n*ߜ� x���ic�	eV�	�u�`�#)��wѾl��e���%��F{�xnM��R����5�x�ꙵ� ���"�&���9a�e�H����&�Z	���-{�a���5�y�fyU�lzB������T!��"Gf�שP'��W�����,B- ���+�Y����.��?-��gt��(�0j�sX��u8"=G�нz�Ư�>�WJ^/� ��Ŀ/�+>�aFn����a�go۴$/����9-#�����CV?S�A��7�]#�=�3y������8�5!�9�\��d���?�MB�4<��Bi�R-W�����Q�V�g_�j`�p6�V���m� �z�u��by����j��*3�&�`������o��!cz�:������2����N���x�.�C�& yjz���Z3�-F��a`Ѽ �mEh5{���]�){[I����T��J�S�x�ү���%)"��C��ugM�gzR�ڃ�J#�$Q��leP���!����Pb�ɔ��UK'�<o1��l��Z��p���˴[P�8ӎc��3� �˩S� �ʁh�,|Ts�o0�˭B88FR�M�� �F�bJ�#�ć0���;�7wu4!�j`�6����3RW"���F��d�g�S�[쒗8��@�V�:�bU����ۿ��5>{�m&ˊv'�Q�NW�'���g��jm�r�5�n<S�HBQ�G���<���$R��C9n�:��- ��i���r�|k��v�*Ilcwe,Wc�G������L�U�X���^A~��������&(����Z�k��[[L>eX�5&�p�k9E�\s8^G!= 9�z<4����7�8p�$��o����=���<5 ?�˷��EB��/Q�fJ�O�  �[V��74���}����.�ntt>�2�o��!�G�?,�ʋ�}���h�n������|���/9����
�Qֱnh���C���>��tT>�gj�g�Y���'.��X��IԋUT��߯' $��r����F�1|��B)���"n��ԍ!ن}�`�q�LL�M�G�g��gO~,o�I��"���Ѽ!�geO���h�F�K�}Na(C�(�x�u�֢�Kߚ�t�0����㰣��,%�
|��sQ�=>	J����usu�x�4w�2�E�3������i��	����R'�g߲�����P��/�L.<�0
Ֆ�MLl��m�R%��Õώ{'rpE�N9H���r��u�M0;y�:Y���hO���<]��5_`��F�������q�6�t���������8��MoQBl�ǡ�J����:�ʦ��������և���C��GQ�ؕD�>��Ѣ"	/��V��Xc2L��ۡ�!�q���H��7u�w���ߋ�I�KSU[��\GܸU������K�	#�9�ڌ��IƷ�]�+�x]4B���� q���� }/tTt1���d��`K{%-�1� ��HZ�t������Է5�Ɔ��6�*�O�����0[�vO�\w������fb�7Y���V&�9r���ZxzTS���[[m�BuP�/o��i���9]�k��Y
�YG�_B��g��x��\T��ψ���b�y�F��2�fOc�4RC���!�R�H�nN|��9�N��x1W"�'R�&B�]یa�MS@��f��F�_Ee]�6��㇛�S(��1�aesZ/��K��3�_ʼ��s�]�#�.�זS��RѮ7졏ˀ��WS�,�h���d�i�46��C~��ϼ�U��CV����Hk~Ӕث���2��ԟP�$Y�Pb3!J�:���e�J����GUY�{�e;JH](=�����"
wx�������k�2�؅-�V ��ֺ�tt�����Ө����o��?_�y�k�#<���,jB�&�ч|�L�f������:&�]�fn:z[�^z�X�Ƞ܋)N{�zćD%��;���hn��m)�oSf�D���s^C�r�=;=�_3��SQ6�!?��jtC�a�	�Si?���W�E��c�g���x�o��K�7��IF�Շ�ERVA�� ����|e���[����}`�'x��m��]j7��/�9>�[���BU�l8zNn+O�Z�:�pa�r�(�U�e�\��l�G�䭫ȥRu �߭H���x�e���C�=�*HޕZ>}(�z��N��8jV4ˇ�g#K�u�߰��|�.��8A��9��D(���}�a�W⤩kn-��j\�[�������oBw|]�-H;��gw٪t�yr�C�*��ܐy"ß��?��k��H/��{k�-Ǹ���X�|�m�g{�y|��o�lO�β��g�_�%;*�%L�q\��>-ǁ�'�H��ؘ���E_��Y��W1�����h�^�Bp�"���3�����i��^j6C�UA�}��z���ھ5�����ǫ����CҖ����e�h�:�>
�?���+uI�<[��.ݩCfKC
�-hq*��h���6��Di'MLlk��.�!x���-D�0�������As���/V(��e�-5Lhs���߲u��j�W�Z������93;a&sx��|
�~��gO�����}\�?n�ƍ�"�W]�X9'�u����M4g�TaV�1���5��8��V��5b�p�� q�\z�ŀ}Q*�εh)$���(#<��	�zJ9��������G�!�-�N^>�^�4IJ
���^~A���{���ej>��X$w���g�U�k�'pO����Sr�էL(	йyA;��5�#a:R�5�K�P�7m\	s|an��=��u$(i�}@s�@WqMõ�o7I�bm���Rd~_r/@��H�2/l:�
�y�}�����t���َ�E�k���#�w��2���<d��v�y`?�Ps�V�JN���@��N4�c������'���ݐ#�~��%� �.�~.`9�Y{TkE%"���ŀǇ�H ��n?`Od�>����a#<0�V����}��>N���w�<��2V6��)�Ќ+�;��{�
��lZE���b%������r���eIV6�n:�%���S���]L���:�������G�A��ߛ��T����>x���c�dpR�\����Қy -hpTv�:]�1�Q�����sa�%��~��O�1�bھ���tP���)�'�괃��y��X
����>H�O�]���bf�vdf����+�uoRvX_0�Sk�,!Xr���U���p��G?_iKB����D�}�����)�1�(�S�[W%]����?5�[휺��&��KW�+�bqoJ	�7�t>�0�W�u����I�1�y���,_�q�`��Ь�|�B1n�cޏM#ȼ]�ƹz[�	��-ֻ�b�n8u���nh���\�f��lC͂�{6�rĊ̀�c���8;eT+��z��^^eQb,����v?���Wb��*$������!�V��}��"r�_BQ���_����x��EQ:���r��! '�;���Q.}��~db&����p��e��5NŇ�4�&�3 �D5S�F�á�'�z�[�i�N����à^P1�s\�H���J���bw�Ą,W��RK��sV^���b�矇�[ኙ�eC�SUh`��*�&� rfa�ϣށ¥���Sd9�^�wm��[�I����x�C3,�ݪa�2��5����$���>��j���-XӦ�1� ����r;=) V����Wx���ċ��i�R����_I;<~i5h�)�4;�s�#b�5���l��1u{�倱)�㔸��Y,;b�ut��������.�KyB���XI���A��z%-@�z�B��ߔ�@����
����S�t.0+dZ����d�hi�r��.c��4��h����*�<E�������]�^�1Հ %Ƌ;R�NZj���1@�[C�*�E60%l+d2R+Ә�W����[�}�Vj 	�B��|�Э��rX�/�=K��0�6x4��M]���@Y�P�(`����1E���z#�
OZ`'_��CD6��;�*���b�$e�U�g�*)��~+|�F�L��co��Ojdr����S�����pb��=d1W��ұ���J<D���Y�$$���8�f�X��m���Y{IAޝ���'�7�g�W�F9B�SZ)+�T��E�ﰧ˳J�fTA��ڨhKe�K�N�P�^���Q|<z��������(45�)�gH_D��cD�+�L� �}�m�O�S��D{�'�L#�l��];@����x�k��9�F�gJ���w{�o�D0q�"�{K����`����V�K�[�k�}xo���>�tj%?� ����
s��ҧ���NL���վ�G_��q|}k�+cJVv:��ch���;/���6����u�����fP���}eȣk'	��˾�@�l��'נk����غv��ފ������C���	�1�c�\�A��5ÕJ=C�^|�g^	}5�a�V	'_8�n7�Xz���n���π�}i�7	.g�:O�:�ԥ
�y�e��7�V�^��{#� ��a��6,�U'�+k��٥3��F��H��]�ؓ`�܊لm���h���r����Z��ME�QQ�^��$��CŸ0��ڗy ���0�J�}\(�~ϿMЙ��'{�d<ncc�"|y"��e\F�M���l��`m�!�Q��C�΀:D �Xer�\9����wd����i�c� �g#Ki�#p#'��s��B��;�69iw��̆4���Ԃ>n.M��e���mݑ����f2r>"N�5⒄�{����S����	�BI����� )�u���`  |��U�&��2ێ?	 I�B�����V�[=3y�������!�
����؞�@�)��LTP��Hˋl�9\5��}N�>:,���7���"��h(�v�<����	��1N���`�Vd|Ɂ�T�����U�$^,_����4E�$�8��A)&_�w��y�W�Ҝ�%C�p�rc���l�
���Bw��G���*݌O@��G�����+a4�J{�L�g+ďx2R��Mh?5�si�i�������`�L��Ț���jn)��\���^�K���,,p�N9�sq��Ya�!tE�Z����o\O�5�)��0/E?�u��J+�Uk�0PB�}���҈�Wu9Y��­�кT'n�H��x.�o-ʎ7v�B�h����d=�F�-�<�/��?̌��Pf�s�����j{M) `����b�[��2����s�ށO��vqR�h����tN��K��D.�V���s�9�
��j�z0ϴc:_����o�`��ꇢ?!�b\7u��{��H��oz��rWz	Wح:C���C��}��&I(�U�����e��b2�|;���F�]�E�. �S |��r�!q�$e3�3VZ* �TB �c�nm�����Y?�Q�Ro����֫PjSu�?���M���R/�m�F��]�Ɖ��m��U:���lkה���W�$���,?~�������{�Z
��a(��=琒+1��� v��)(��[YӴ��a	_�RkC{bc�/�徵 �a�0 ���h]؄�to�h|~�6P�� '�Kl!��uxu�9��ZoY�ԍaW��{W�m�u���E0�&����=_���.U'�$j�������*=��X��k�]���_[E�tB�7(�n�јP~�_�ې5�k�8n/8%N:Lg�C<�^������5����jy�p�D�m�h�yq���A>鴰�M��i͎�N[ ��`�-k](Z�7�@z��S{g�s/���Ң'�F��Z���vǱ򚑫�
��5��H���m�o\����T��鱮ă`m�f�2�F,��G�S�I�{F9 �M��Q{e	`f��6g��6&�<%��>�R�v���Jen���4v�r��
��0 ���н���F9�E4$���<�W��	��ۆ�ѿ58@h���������q�p5��{�U%Է�M��.�TL�b�~�+!�dD�4{�����A�G����2鬆�K0��_�Xl+m.qB��\ 	��h�H�Ў��"���_}�L?�f�YHY2�m�Wo�����i�Vê���ȑ�&��ƨq�u!S�s%@| '�[����ӬW��tZ�R�D�j�r���۶�ks(��̤��'v��3)�TY���3����h��T�B� 9�V'�*���*���)�x���#���;w�wB��R���z�z-E٤�ԍ�ݭ"���e�D	lo����5��5��Uq�S9(b'J0Uk:02�rD��=?֚CnS�H���8���;h��v#��I���4ɝ;I$a������M�l������H%�:,S���E:�j�W C=���礈���a&+'e>G�Z�ݧx�,ӭs�4&��ݤ�cz���o�f�}:��{�����9���"@���=��Br��C_7I��z ,=N�<C���u�~�&��Q��n�����sZ�����:/ѝ�U
	�֯}M6[�j흜`� 8\k�pD#��ۅ
�ɬ��_Ġ0���8��iQp"�	���=-)�_0n��n%��9Z��Maa�y��~&�.���`&)S�y�m�x�"s� K�t�7�������P��;�ϭQX���z����7P�/�E讨��!}Sj|>(P��B��|fB��)�Rx�O�+�	�^�0���L�����b��~��":Щc�!���2P�'yR�\���$MH��`r>�V���ޖ�Y��)veC�����6,&�t0&P"<��C�|nvo�Xq�P3.�&5��MR�(G�?5o���OemZ��: �����<�RZ��cܶIUD"�B�u�g�k2�9 ���Q�{mlx���Y*a�J`�0��G�Ql��]s���洷��U�P<�⑇ۅ��i�I��e��{��eoҞ� ���H7��<?�sό���Wn'0F�� ݉��_�(��F7eHQ����R.��ķQ����%
T��g.�<�M�[���uƟ)�D��"71�<�.��9��:�;� �G��Mz�	O�����7���)bK���5�5]�Dp3����
���D��w��n��X4D��|
^����>d�Ak)6�70^_�\����3/�Xeo��Nf��^ڄl�Ƨ�^Y��~�����C����q��ëi�O,%i��ovj�&�\����g�뻛�w�^�vѓ�;&Ӌl�^���8zH͈z����d5�P��'����K!�S�.�]�O�r?���Y��������>�Ǵ}����9��Cp���lh��~Y�j#N�IN�������l�RXRC wc���J+n��iV7��@5Q�O��lX����E��2��1>�6-*s����ʺ�{���rlr����&|���� &�/?m�#̵�z���P\�G�<�52�v^�cjz5�w�)l�\��+w�I)�Ti�����.���r��{W�-т���蝹�w#����n�t�P��`b����'M^qn3k�>B��2���������ZӦ&,t{		ktB+��	ޛ@(0��(��TZ��o3g�C����N�3ib.�a�a_y�=1Gl�iʻd�YӨ�J�����h8M�G�~��Vю8g?����EW#OSP옋���5S�WߊZ�t�ӌW��t]MZ��㪘R��Aә�~���ݫX%�6��5YW��M�!�3�m�>�6���l�T��P�ի~�f��w��3���Dh0��\��y��y2�_P37t�'��׺G�y����f��łd�t���
@�`M���a�o;h��U���n�$�
k���}.�'О�I�S]G���b��_Siiu�yQX���ꔘ��c&�\����J��s��|e���͍��� =���n1���d�Y�Ɲy� V���h��1��xp��{Kd��XoW�#|�1�:�fH���̕��gN�k/���b��*?�~r�ע;A��e�y��6���(�8�|�y6.Nv_a�)[�6��X��Z���#*Wг����_:�А���j2�,�/�~�7�_�M����嬙'�W�C:VpTDN-�	��Qjذ�>��"�f��@Q���3���o���8����ߎ�c���8�sd|v�ٷ"pp�Sۜκ>�y�J%r��2��X��AT>��%P�e8���ó�c;V�I9WS�Wa��_�R%��Ŗ!Sޑ�E�D�����Μ(`xt���A���B@[��l��S�ek�e��(ׄ#�D�����%&O�4��8z�Je�C������0�pGT���@T��M�Hļ�ń�����P$̿M�_�" �0;����/h��"��.K70��BL|�^��.�1�G��c��].N2f�����`�5�}w�(К�`�zz����
Mc�-��8�O��2��0L�oT%�:8��>�g��p��[hum�DN]l�b@�ij��lD�/PvvO	/�b:&���Q~�ӊ�*iaO?�@�~�@�t�k^�o1{{�O��my�5b6�kpM7��Q�x屧9�ƀD��M	:Z��m|�#R���<`�/�!�~cBJ���X��ԯ��q-��K��,zA��:Tp�@�c;ɾjPw`���ן�%C���|@gY�J�q�$�������h���0�.����c=��9&�lZK�5����[KQ�j�Y 6����gCl��F������H�wQ?�|������Z��Bݙ�	(f$g����Pp�镠���<��IK�p2�@,^���yԩ�P�K����?��a;V��{k7���X�kAu�rƳaB�y�L,=�	)�������G�j�3竘֖Z|=��e70�_��c�+�it����F0��%	���q��'�g�3����T�a��;HA�Aj�,��Տ)0�г��h;���T��Wr������z��>^vm�`I�wU�["O�.=p�!�i�[��H>�)Ӯ+x-�Ě��LL���a��M;�xT���G0���W��j$�i%8�b���h%����rQ;��0 ��d/�:ŋ���=�S�������Wy��#�Ӕ9���P�����n�U��d��я��f��MQ���i�����R����j�Mq�d�؋9�?T��� ��M7���!�8���e����rV�bZ�W�2؃xȗK�ں�p~�8X�ﭫ0�A�vAD��ق��JVt�h��ϒ�z4��ˣH)} ��$d���J�~q�Y)0�SX�s<�q��Mݩמ{[����Q�@�=�
�;�v�|4�A˒o��o}�w0�/R���]'�����$�c�r�zNԖ*5:Zq�|�&�;�Ԍ8W'ܐ��aM�G�#�"�xŇ�Mi�Z�	��> 9��+e��.����t�bc����P�tQ�z T�ԯ�.g����7Mtb{V�ŕ���KbŶqp����ׅ+5L�n���X}�W�����G�r�Z��p��#�b�&��r���M�)D$3ӣ������y��1�l�B��`L{�Ɯ)I�� �t���T��ű�=�d�։�2'TMr���8~j�^O�@����q&z�Ǿ S}��i2|)t}xy��w�?$��!��S����l\l�~rN����d��'���(�_����z��%馺�a�4i,]��x��[<b�gD�ɼÄ�<O++�X��u.�\��_עjx1B ̛���,9t�
n���H/㤅
e5����@��� ��ݍuH��䊛$[�i�+��V����nLu����k�?TF{���r�as���I��2�-�(q�E���~-"�n�����&�iZ���q��HZ�.ߓe�(c&zlZzq��ɛ�ԗu�m���5@DX JѠD#������;�~����~�->���a�/�G"͙��m��<\f��������)W���`���0��8'�idЈ�Lj�����|j{zkѬt�39�5/{��xn���FU�k~����}�E�����Ws�}���0w������x������Y%g��k��(��iBL�Â'vy����������$>�VX���}�
(p �;$�^�a<	u�9[A��f��lKX�&�x������}�"��s����4�}�4ڱZ��n���	�jl�/��U�뒍��h�#�Q���Yi�m���o�'�|�r�8X'O��-�jqFT^KWm~�uj��nɜp�_>� ���9�m��m�c��2�I�È�>�-y�g,yEY��T���]q�PAo�!���?-2B��3	c����M��S8�Y�"�m ������Ƅ �iQ�k� ��7�w\A���盳�2����		@�|�FY���W�i[(�џ� H f߬�t>7�������~�:���������;1>ɿ���1܆#��E���|��H͝���\��n�3*"�b��pk���r�l4���;�N����-�ݳY��DRðɔv3�D���!ѱ��%Z�7�D�)�����e;��C�H/c����:Vju�qK�n�;��u������k���5�l����e�=�W��QD�՜�7P);����}������}j=�͛L�ѷ�:�'͌L�a�&�a�u.O�����l����'��F�>T�?��)�-p�`a�'.��F�=@f�p��|�&��%Ĕ�a�6�Z7�{�8����f�"����Ȝ'
���n�����kn�N���E`�0ye�T�G�\C����/����`�)� FT���c6	����ۭ��V�q,w��o�,O=U��
v���Sjꭩ}0d�l�ǻ}{Kv��ګ�煛;��OMc����3m�?����N�lUu]�p\���l�������-`D"�_n��R,�O6�˩����-�bF��3_ֿ�1u �_K��d�\ _>��X�QB� _&o��1Ұ߿�|T]6�$9cs����dg�����W��u@!9�rsвz����{Z�B��"��5��\�p*�kA�}����w�FJZ�j�xW��A.E4ƶ* �m���Б���ů��&���׷��fU߉E,4 L&np����<�k2��d��%��1x�O�����06���cj�ߑ-����1��,˺���i�[�j+��
�7<=A�%n��u�~�+���I`a�@O;t�ګ�������j�kS��QlJ9W���u�L����m)-խ��z���k_��^i�޽F���t�٢F�P���D҈"�-�7�<֎8C�Y��?M�E�p>\��W�( �_(x�85��3�xU+:(+�����a�?o�^���tU���k�?Y�V#d����k��s���F����s�h�Ş}@���a���J�|���ٛ��h�^�C�:��ϼ�j���6ɕ�Y��*��l�ȅHLm}��(vqlP�H�W��k�0Ū.ߔ��I�C�S���/9�<�Tz>�$�1rF�O6�q����{���gwSȴ�M�ˏ��Q��~�T���Q�\O�n_�b���v�� =�լV���:lN��K�
�쉭�`B)MGC�D�tD���tQrb������7�Y
�e�� 䣰��h�d_��VY�����`1k_;�N��S��ɚ��Z�� ����o��)�	�Ɏ�EF&o֨�!����9յKn�B`1N�nY��H��U��T�k������tv����$j��z�_Lq<Yn��2�����;�V`�z�=]R�����}�Y�ӵ<1�a�NU`�żz������X	KN� ;3�̨�Y��<�Sə׼��p�}3��b�U�����Ve����_r��̮,���e6泶��q)F)�b�G��R1�� Kc�eէà}��x�������#�;��z�7�l���9��o��+5�'�S�F����we��4ĝ���D��8w�<�}}�Vf̎=����x��"�a#-��]�Ж���M���_R\���^�8O��B�&	�$�Q�x�5�'��o��z`h漠�Q2� �?��Rω��.E�+x�n���^�j�1O�mz^���/�ܞ�*
!-Ԁɛ`�����9Z��5^�ǪAS��T��� n/�G����b{i&�z��٣镥�;MFW�q��9��%���s)�
���H8)v�rE.�q���T�*B�hon��;! �nA<Vg�1N/��众(�`&
�{�q@�r�����|�Ӓgb�[��Wd[�@�ׅ{L�@v&���������D�>^������e̊��>]6����a}@a�̎.PͥP+K�O��xz�9���T�y���⪈�H��֬����B�O<J/�)j)�@2�0y��~	��� ��e�7eB&��d���`���!�$LQ ��	Xr�
^|��gP�5�����e\Q��_J�Џ��OAxŠ�wB$�Jͽ��Tx����X_��ؐ |[�~��
c޹g|<�!j2@#���}��iYܾv�S�_z�����|���W�d���"R��ׯ��D���@�&5[4(vۻ>`�<@��W`���#�cs�#e�1����i[!����qm�[�8t��\[}򯆬�D�Zj]���G��jb����oG�p�*��6pXt�/#�l��΁8�w�Mg��6\p9m�n��X$�f��,F^���I��J��۞;�9B ����ӦN�e���*ʏ�̷���:qQ ����|u�>��o���p���v*�"��J�qco(��;y��}�ih�: 'S���惯Bck��w��/i�K+����&Q&��RUl�4�w��WA���$P8��h�%v�T�}o���J��șa#�Z��$��`�����r�#��v�)k�w�Y@egvh黫/,��ʊ'<	Sh�.u���"^���"��a��	]�9����SC'7Y�&(z)�*������Rә���W����,y�K�Z>x��%�R �-��qd8�H���ns�4�V�V�t�a��s��c�Òi���<�xfY��g9ϔ+ o}����R���G�`�~�͘���Y�u��p�e�z�ޅ����a�z��<�/Onr�f�.?̟̋�.�2""�fK�����"�N��d�&E$���z��i+ ���w��e���_�@�Q��"��vi1�J{-�׭��7jY�Æ���kK�h�@r-�H�`���;�AFL��w��6����vZ@/�꜐ҕ�A��2���*/e�(����&�fd4�H�����&�Z�iv��@n=�j��K��Z��$-�J�K����`=�&-йƛ�ى�~�w)+D��꺚q���f'h�����)�W����h����]���soN�e����Q��P���u����������우�݄�
�vC��L_Rpkb����F�BDL�"�\=)�a����)a�,��!�ٵ��N�)-������H΅TC�Է�ݴ�O+oo	:yd]f�������5^������{+O��X�n~9�T��Y�Τc�(�O�1^NC�U�EoRDf/i�p�D�̓���� A��)��a?��v��7Q����|~gϚ����B��qQw?���>��8fZ�V�O^ETq�L U�U�G�v���P���fP��-k�m�`���Nl�<;B?�4j��0�U<8���h�:<����rl\@�0#m��� �(���W�r1��%�E�gP[�I� �=I�igݸ�U��F@�DM|�WR@Ȯ7GJ��fkS
��6�%�f��<�XS-v� �u1�[Ϛa�k��CW��b��7!��s��h��n�zAM2�	����Q�F�q9���CKx1~oP��Θ�~+ۡq�E4�~�������,�����#X��6�g�Z�h@�pC���8��D�3��x*h��C�-�;�R����^ �GT�m�y	iV�3�%Y0�½R�]�>ࢎ�u+I��r�g�r��WGe���$�h�c/(��S��Y-���ע�L"S��|&h;���	
�Q���X��.����l:Ц}���wl��J���@�W� ��T0��l����+�d�©��-�ԙ�%0�ltX�?뎨�u��c�:R��rNH��E�٧߆������ْ�Y~�Q6�����]?�K��Ƌ��l�(������u^����l�K�!��2c�#���5[ïܻ��P�Ku�Ǵ&DY(%�Dh�|xn �b�9Pm�R����9�<���h-���2����-B1Ͷ��Q#d�'���5�q������a�\F��+��v�\�
���m���Ț�>���\ξI��G��Y:Qv�!�X��p��7\�ȏS�^��G�e�{�����b��S�17����R$�i��H��˽!^f�e�K�i+;v��n\���y���	!T�FL���o��qy��m~���aq����g�7��w,N���)�p�����W��%�
is��$�ZQ�
5���-�V���y��M�̦Lj@�$�P�qp/.WF~���) �����N���k�r�o^��b���Խ�vj��E��UsN������&Xeћ�K�-�����6r?:�5��?�:��D��T��PuX9���1~ɒ�";�(|���l�E��a��9LY"���FG$�7[esE�*����Kyk��D~
��yO�,���y��v(���g:���"��m�?X���`�@v\Vը�l$q�O�?�q�o����+^�C���3�KWX�c���u���5����{z���s��
[1vn�~g{f������[��_��;�$�-|9��I�)�Z���>����$��9�F�Gt.�u8����Taڷ߷΃��7��WQlå8�/i\�_��{s���lc���eYg&#��8L>���<z_�Y*�|r��z�I���}()�\�Χ����ڏ@�FمGKy�2A�	~�4%!���]w�YV,r�?�u��N�4s�t`m�-�[yޤ�z5{�I���%=�1�IV��m������w�!��Gj$��/N>C����=M�E��hg��H$DI\O͉��G�����`�K
9����aW�~փ��d#��@z�s �!���8M�ӟJ���K#�����?�#_���U)��(q-ূ��-�Z��GÆ_C��h]�6O�A��jLɈ���w \{�
e�cƮ�nK�In+92CVe����8�I�hoD�U�J[U����,����Hop� ��d�$��8�0,3NῸJ�$軞�.������ra���Ӡ�2a&�����x�^N���r���<݈��&{wI�d�+��]#�W[7u�Hߧ������{�A��,�]؛�:D;�2Nkn���n���?�k"����НO�۳շf0%%\EO=�m��3���9J���'B��^��@�hZ:��f1B�ҵ����d��U�H᳞�`��ZH�oa�S��v�K��54f%B�JX1u���T�s>!_�*&����"�V������R����5Έ_.��o0-��^���I���*O�R���<Z��'F�d6���jyT��K�6��Y�R�B�6�UhQ��7�9��?�ն8����*E3R�(}��#���W�. VT���@�X�?9�LJ�/6�8?E�|^���LJ��d�[��m��;A�ahv�F��Vw��?�	O1���ja��-oq�̅P ���������e���W�Y�����3?����8��H8��Σyݨ:@5Z]��I�5Λ�Ou ��ZUo�_a5g����˹�6Ԇ���O�h�sVh@?�G֋x���,	#�_���Vġ��Y��p?�$x�UĖ��ZWa�)�IE�Ƹyq��}�h� .��0g�j��oK��m���D��;��)�������d�8�&0�5�C��y�3�o�F����Qȍ�j����@�s�䈓�C�eV��%4&���=n�ԍ�4��Qg�5I�t|�һ�]�ѯ���:�0����&:��ѩ�.>��*���t���陎&��7�.E��5��6�r�@����H8��U}������2
���t�	��������7"��:��<N���x��F�j�7X�ٽ��]��IS�C=����	�6�j;���(���R�`<�݇#
�44*�%;e���1<\e��q�&���f�Ȇ���_�7��ً	a6ڒ�f*��mT>��%����B33�|:���������L����R��^v揶�=��1�W��2kO�����&��k,�@-,��ơ���r�+���L"r-��DvEi�[�,���۾gߚ�K�.���
��$�iK�p{�Ȓ0Co�B��Z~2CE:�g�<0��ә^@�� �:R�Q�2:��P�:W�0�`��g��U%}���*�X�+��ב�])ǍP5�o8�!x�*_�G$�U:�,i`� �ѬH���SeX�t^�_�~�T�7:_r��$ċ%2�I l�2�T����ֵ�:<�x��^>���c�ޅ� �K�����C�����1<�~`kY4ؼ�sx:��|�ݒ�%iNZ��I������D��bl�F��q�צ�tݱ�m�)����qg��9Ͷ?G6N7
V͙{8ޒ�$�-�VC�s�4DM�7$f��H!6�V�Je�	�C#��+�#�%�;��5:����?8R���`4ll��������&}�gN�>!�5��?P^kՓ?�#O��˟�4xh�~9�4p���e����#�o��I�����)N	9ݨa����E�������
"l�EYuS.EB����0 �l=W+�I����I�P�a�"Uj����
z?�mtu���9,�-a��H��m�4��j��n�Hw��P�*����׫���� ����J�͐�5�C�3���pN�o��_D�oچ�E�Ni�S���M�����6���~��F����/��TW�H�UZJ=���!�h�f���쏅 ����,�q����iѐ���B�_���߮T.�>����78O�O^����0�G^�:�_67�����$8��<Ó=ߍ1�R� �����cK�"� O˖9>��c?e�԰��Q�e:r1�%"f�Xʳ��kA��"���i�G���	����:�4R=��!	؇�@�8���o!����s֢*�
�W´w�rã0�7P��t��J_��$p������V�#�Z����-���ݰ�h���ݷ-=Jv�7EP�4�/R����޵�����v)��q�y�$X���s*�v�s�Vŀ�҃4�^e�y�W�I7k\��'	��[�ŵii�V��l�vHӶ�����W]k�����7%�����?�gxf2ّ[��k��a��<�誵: ��d���*Z��֒1ݐf�k���b���1�g}a�I�8"OL@��������{��Ni�&L7D�#UIϸ�b$6T�X�I,��󮋋=Q�Q��
U`���:��̛)LX\��H��ۃ8�L|>��Ps}
:+P-|��5�&�xRX����_�ѐ�����!�x�zU5}n΂ ��ϰ�BZ,�~�K���{.l�����r������P��F5��)Y��K#(R�&A���`6BJ�J�[ev�|!�%X�����Ζ�_�I����ph���E����ݽj����bH@=O��`���\Dx�R�tI�inϟ��x�712�*�Kr8����ef���}�A�����1���*�͙F�_�r��`Q�������$S�<�t���\!��[���>5'Y�jWH�^&����[�����0�����f
�;�Kcnr�E[Pu��������v���	��
�����_CSUD��R��!��a�����1����ͤ��We0�)�����pҁo(��-Y�,| ʈp���>�R�oG՜cڳ�R�K���4z8,Zh=�L�4R��B���7z$�Ǟ�=��k9A����i�/����Bv�\�/�'����u'��-L\6l��B�,�ж`)%�������:�Y��ВwB�o�H���z�ᦤoE�h�^I"%�	�6��f��I�mq.f���<����%�	$�����
X��=�&f�����=�<��៊M眕�����.�(�:+md{��U *k'P��-	�J%2�{"-����q���Z��>͠k�Т��=�p��#@3Or����d��Vï�$b�W`���2J{�[q�"" ����K��%R)�G)���dd�(��1����y̰��*��)t�	�5~�Hd�>���"�����:��ꔵ��K3��g~�P�$�3���,��
��Tt��q�	,C�x<�3��]*��XR�l>�(L���'��u��;,��pnzi�r+薎����isQ&�?�)j�@�
	��Z�2�aI��t��r����`1��N�ѣ&�b��VB�F^�6Tn����Kto/�yf�|���,{�$�euqFs�T͡�錝Ð�.�r�W�7q���zN�a"܄j�־��ĥ�h��'�_I����(��:�1�,[`شJ�۴РS�s����]�
�zi���	D,c�Uf����-�I�o_��F���ו����#>����D�X���&�#Y��q�}D��q�he�T9��#4!o-�RnL\�	��]�PP 9���p�p�q���w�I�c2m�n�����$B(D��0B�*b�9we�Pͧ}�0��N����Im%��cc��jT�f�q�vZK�vq ���-DK����4�6R�?�e�e#CT�|�� 0p|;�w.�Pl=N�	2���12�Upqz��Q6����BE�t칐��u��P�k�x����W��7��^.����Q���:y%�ލ/�+^T>����g*ׂMM�E����4^|�C��'��?ά�RTl���9h�#���3G��<2�G��������A�%���bR!���G�J���>��G��/�Ǹ���\Șr��8��6�����#�t%���*�cDO�#�M�f�9`:��)���p
��C�??�U�@7W��j(,P�S��B �3���:�4���5���>�#,����GIUЃc[W��a�)�V�
�'̤՟����9A�T3��Xv���mѢ����m���,x䲐Ly6	�yO>�� ���B��W)�@:�P\%��a�+Fv���m`2YyfT��+ߛ�1�
�u׀B��/�Ӝ
 b�G�Ģ5�+u���t���o��!��g:�0l�-dX��Ҹ����2p�H�l$��ls��$X�p��e?"@�Mm�^�,�z�4��r �s��vd�[�mN����I���4; �ȳ��j�<ɣk�����0�И�(10�O�l�Fg*ES��]@�o�%���=�t�XuH�P� c"���Oy�-�Lh�6�Z��g
C���<SqB��n�`�j���A�Lslx֋SdUeԟ��+u�h#�xe=����6[�p���WnV�i��=�,�4���'H��!��!<�@~GSr�iME��m7\���x H�.�kR�sxKf��Y�Wq�����P	�׫h����<�5:N����{�F��>_ox���93,N�2�NlcV#���i�ɴ�:g*sh�{���� ��#�De���c�6����,�ZK�b���x7mי��!��U�Ȣ����PDCX a�j�$��&��Z�'��.��C[�=�ɻM� �<D<�A��v���7��Z�Hjh4���z[24M^0��o��<�Pe�@�%'�-�@�֜�ȡ �*�Γ�߀��liXѬ2��`���=[��S{��9��ɂ�Ic��b�U�@�t���$É�وW<9�]V磃O�K�J���mfZ��'�����]";�2�:h<է�j�x�d�, k"8ݸ��-��p܃]��������/EpfsB�Z� ��^8]E�	:[��]7'�\f�3��c�*䖓��{�㧈�j�	�C1X�Y��KTG�U��/�]PEat�QE��w(C@�Y!�@�[�9>,��:��O������z� ,���ٞS%K#:��H��M�瀸�0�\$���Zw�>��a�j�uA�t�k��!��vX/��^+��O��h�SL9@��D\�ٜ�/��k8�r(�1)RI��*����4����N��S�%�F�M�TN������Ү����PDt!�p����ܝ^?P�!&>�g=��_¡:D8��<�7��QNq��=�/�*tU���"�����ĵ�Y��6�VUDIdӟ�0�@��H��P!��@O�(Y�Z��s��3Mg ��V�t��fڌ���������$fc�JP�wZ���������`�q����h�^�$acKx���
�O�*~���MFC�!T뭸P�j�pu����:l^���x���: R����C�h'p+�ar�f_��d���,�}�N7������\��zHa��K��T���a�����a�EcG�o_��N�X0/�V�Ǻ�9�)�o���Ꜳ���\+�?so<m��G�C|H��Tj��ȋݔ�O����IFI(	����&}(�h\kI理fe\m�x���Ws�D#-�z�`���iYe����	�|��b�G�5�ҟF(J�)k<~��N^�@��0}��N�1}."xh��Nr��՗r��jՉr�)bo��+�,��@@� �Wn@*��7TF*�Z����{݅�!�9#dxJ�Ʀ�e$��NF��N��2�H���M'� ��N⟧g������h#���S��jn��Ss��"��ɦ�(�"��\6%۴1���5 /hx��C���9[��3B����p���Ň��B�pwYͷ�18a*;,���Ī�$���t�u��������X ;P�.$㧌}��K6|�y�hC�b���1��x��z�ޣj���^C���˞3Ɗ��L��[�|c�އ��Si�d��K�?�pꞾ��b��?=�ðsS�����L�<;�S�P��#J�C���/��ԕ(��Ѻ��>�L��ꍠ35�n�(�� �Xq;3D;��ec���T)�m�/.	ݵ���"��d���@eX���/�wy㿷O�{i��}��>��zi��Wj���vM&
Y��P�so���]	�m�:d*���$q�ޅ��:�h�ǐu[�W��L�E�Pk�e4��@�i剴Q���4���E Q��ע^�����
U+&��y��5�v3��#p�#p�����T�@o5Xi5�����a�洑�%�8�I�_� �+�D��d	�@�$��U�m�dC��_D!톊���B^x	SH���)�s�I�7wVχ�޶P(<^��W��n��A<��S|�8�/�-�gt	�$	�IpӮX��O��R��>}���Ry{s����9ζV��b�҇�����j�o��+�W�k{��M��Q���������b�<�O�.u��V�R�(��̥�+i3�֙3��Jjz�&�Ρ#@p����{����.�-��8Ӛ����.<w3��+�=�+�W
��M��T���
'����_�<�zj'���Ҕ���	���B�A�Se�y�M(�h�5��*//;�C�6<���ţkخZ���U�$�����g�� ���{|<���?�;
�����HR�gmR1��[�Œ��kZ�>վ�as(W���Q�r3�K zq����#/�#G�񇳺���X�0eB��� `�͑�Z	.��'�ƚ�,�i�y�*g�9�i����/w�)5�1UI���X�s�(9&��q��4�V��HJ˻�.%{�q�3��Y� 5
����88:�m�{{A��]ۜ�#T[��4�*�/��h���y�o$�hĖ��I�r�O.���QM>h�b�;|�=�'��>E��˶'BK�ďd�='���F*��|��������h5}�3S\{fEm�l�lߺr�B"��A��k�9؛{ףj��TK��󐿓���P�:�*,y��_�����c�	��(H1_���aK��e�$F��?ZԆ)R/���ȭ�6#�rE�v�� A�����cu��I9MQ$m��������';��1���X2N%���ab�%`�w�M�	lz	�2�-��������8($K�`��b�ګ$�����4�T�u�X����\Ĳ��0��3�:�l�L���@kv-L�VOi�9����+�TK����sNVIM�e�jn�9�dmk�MzJK zc�Ql�qbm�ҴA9r:6�q��a�3�׹"|�F^��]Ճc$�=�UH���.�9sѝdj������Cg��n����ų���t �H�ʘNT0�V�h3�*$Ik��i��<�F��S�0ָ����i�i�Z��竁ܜRT���p��k�fԪ�B�5k�0�8G����S2����
韫�?HF{˭k��O���>G��S����X�p~��W�Z���$�+�ӡ�|�� ��k�\<  m/����NjhF�D���w�* ��[X�U�U��Gd{�
�
�G�����%��&U��o�P�w�+�1h�|lsL��U���$�b'۶��߈@�����9;-�Y'�SM��(dC*��Qx5����TI%����f�ْ=,���6#v�[��ܰԎ-����T	�/4 �����A���_�Ñ@%������cn�Sd�;�P�$n��t���#�n�5�p#�|VfR���9:-��Hɽ����L�@"�WYA��[S&��[N@��A���C	�u�qE�i��
Dwb�߄N�� x�"2�w�}���D���ݻ����O`��5�ǲ�*�\�E�!s�[�"<�?'��L��0r{�\�^�'L���dJ@�X@.�o&�ܞZ<UY��5Q��uNJu���"�ql�r���hj��3���v_�>>K�n������z���C.C<�f<A��"��*m�Bj0)�q�� �`m�9nɄ�Vr��c��Ɯ�mQ,��GKb��%���?�qx�Ut���B��Q�!�T�Y�Aqq�������S�`J�(nY?��|��Su#���y�L��,I�i��ćc~ރ&�7Z.86Ш9�^��2F\7����gk�&�8�݁�A����Ç��������*�|����9��*e����㝶� 5���c�pq�X���@�c�rz'��ZRKK[�k�U��o֨qJo9ޞb!�7����:��Y�h�2Ҍ l��F�b+~B���`���kF��ӂ�]��tMj��HF�)c��bǲvI�ވ�>����x�v)񲢏L1�Au�l��ƬL_�fN"�0̥GG`���U�'�;�1�"/�V:G�ߖT25��n�td��%��������#�̭	�t��G�����b��$�����A1����қ&UR�Y�Z5�g�V�׬ LV2��������d��������Y�/�v X�.�;��,��j-s�K�z֡{�ogK�C�/ä�dNr�j��M/㣂5UQ����"�s3 Ipq�%�m'�w���w'g',������Y�)v����X���h�����W���y{hBT��@�l��5q�?	>�U KV�̕���7�9gkuB��%����2� K��)���^��J��$!�qe�~h~rz̱�e�_��.�E�<��7�I~���}_4�/�|�s0�S�*�Vq� �f*�z�25���i<�����NnV�@��r���� �<���Z>�s�m��X�u��iUJ�u�-4B �����rU���H��UW�!���}9F�j���&�dG�wSj���n�2�%�>�Yߎ`��B���qۋ�2*��޷4���I�D�{}٧�+�z�L���Z��
�����*լ��T�����K+�n������N,��9��ѽ�yyWM+�t�O9��0��U�s�F����,6)�����wvH4&�z�x3hR5���2y�-�I{#$���� e��
BjC~�&�m��7��Sʖ]�0��u����X�4Q��r�<�A���L�������N��3ߤ
���� ��yc6L�v��t�9�f�!���x0q(Ͼ��ɠ&i����>d�P̉�����=+�Wޔ{��B���p
�>M+%J��^������~U�����t�O�"���J�i�N�6���9�\���e�k.zx0�>BJ�O\�--W&a��<G�CXZ%��x��6���;"�^|�L�.2��3_��\~��U�AG=�̄ǫ.�-)f�)����Gr�T����K�w��p��Ī�t�p�ыKc�a��m�M�t��ɓZ @`5�iN��)�#qf�CڀO( ��k�UOM�ФE�N�R?��`�*�_g����5HK���OvkX{*g(���hj�Q��S���z.I�KD-f3�-�p�K���A�1~��@or���kHX�t���4�@�$1�K�V�἞4�5����	gx�t	[�d��l�s|���ImY"!�SH�NSe��yS*e��i<�%A�V
�	��z�D����W�>�t� ��D��T �h��+�s3�J%�-����/UybK평C�[����]�#�KtT�C'�	b�ʘ��e���e�]3�o-��$ʬa:�F��'�	MI���;ǥ�ʉ	�tn�r����F����W�eT�4� n���|�SsT�T`��c����ڷ�1[����@�>{YR�8�܋�.�`m�>��g�����5�5�@3%8C�a�ԙ���f�I7|�Ga�%�)&Ƞ���秩�>w Go����u�!��fS����d���-l���[p�i.n�]������_�Xx"Î7�[�Ѻ\���9� R3�/��AB�!M������D�b���k��E�?�z@�����-�A�������F&�Ս^�}�f��
�u&�{I�X�i��v�D-� @9����[��'��JN���; T9nZ��a2}�,�� �4�e:��2�}UY��/�E�vXD�
T�š���?b��-��b2�XL�Z��,�!�^� @�]��ӧ,{XGW5�
�@�+d��hN�~�λ̓��P �K���z��P���Y�93#бO�V sǃ���fE�ؖPa��,{A�7Č���'�_M@f�|��M�'��qш�=�3�,�-q���WҐ`��J���ì�����$���}L���x���
v�D�H��ƅ�jWp�%��W[�+��^�I���L}��!��A�vi�d�u�[
_ �ޗ�^�m������#��w&�QUv��#���;��z�MU>���tX����D�cq-f <�ײ?�k�_y�&;�e�z�n�� Vmw��$;�]�T�k��2��s�����D-����.�1�Us���v�l�n;Q�'�akT)�]�(��K�ڷ�M��6�\*���AMUp��L��ټ�W ���
C;+���@ۛ�Q�B���G��T�L�dK��Z��u���0H_	��k�Od^|Z��d�p	����/D�DÁo=癋��aOۘ]r�
4j�QɿN�h�C���=�D.@>g*�c&��PJ���Ǣn	Z�+\F�8��ᑰ�h��ׂ���)*�����X�:����Tdw���� ��K�B|,��Ic]�Jp��`w�\o7�D���4� >�V����Jr�1�K&�@�ۤ#ҎA	μ��+����ṙ��|cDyM�H��S��ĉ�{������o����lT�+�����N����6��6������
^OE���wŉ���"/�8*�5D��Ȗ��_B�ۑ��1/s��܆h˴bfͧ$λ�4�C��~�-�W�^��YNj�,H�V8�b�1�szl�p�N@&jH�;�>�)�p���x�Y_�<3\� 2�I���ajx?�r�gى�3�$<�A��q�NF�3ğ+�%�����Q��V.�j��L����wN>�лi�Z<���ena�n�gn�q�dŎ��> 4�ݼ������oRĢ��y��Y��^FǸ����n�р+o��)$X]�ɟ���:d���&���3jF�����	�$.���x�0
�n>��S8��DH8Kt�]TɃ�2{���`S��\'u�1jy/��%��$]�Q�З\�>8�.%�� m�t����R�*;�'����T���!�}}���L�R�+Z��KY�P	�kCy!s���z�:M������I�#����x�\0&��:\i��?6k���;u���:�*�uo'�R'�jjJw�@Dox%���]�k�N�)q{	�ᚒ7����J���mR��/�嗿}�]�m`��j�f�GU������P�����Be��!Y��Z*��q�JH�c*�S�^�6I�3,��	ĕ�ӗ�RD���Pjס��3��&-�04���*� ���`�^���	�5�g0�*dd$�-��dvF7���O�p�Y�� ���2z���0U���s��P�-�5��Åv�tu�No��X 	�td���6�熕e��^Y����ԟl�jg�R��:��i��َ����I�Pce�U�7��j�kC�/C�:3d �F�z�0�E��������S���'�
-w0:=3<״%�/��l���t�+r��ȹWm�틊Pt��i}�#�pA�?X�B��Ay߁\��:巠r�bkK�����`#�&�㾁�O���6o�fo��j��Þ�0,�cҼ"���7?��)q`B�����hю;Z���ZDe3/~,��ӭ��7ߓ�"O�8��D6퇔"0_u(��`�Wo�ղ��!�7����[���+����.��i��b�Q��\����2TU���A���K")L
����]�t��[Cx�ΰ�ӝD�<��l�%-�#�Xf�cz1剌K�4�e/K�ACG�N�����x��D	�$��
�x4�T�T�-.����}����y)k7�y$y��hc�����{W��JA��L2ߍ�O%��b�=�ހ��A�r��nuzT�%5�>Wu��\j2��hO��*6@�p��?\����#,���$a
3F��<Avޭ�>?f�=��w^a�C۴E"ƙ�vfH`��N��c�e��`�;��S���l�]?��}�;���&k5�Wh���;�Xf㶜f����p!G�`/�sr�`G�!wx����:n5m>(oE0�{�"R�k� �4�-jm��`��B_�<n>��(�4r�B�Zz��C� �E:����o��!��ުm.�x��T�؏�߄�X' N�E���ᛜ��c։��_e�)}��Q�f�%�ɉzP�1M�/�������H�^�U4�bA-���gm|���ؽ�`�I�3y����S�.dBł�s��3&*��_��b��$t���̄�/�������'*2�����b)�!���æ)&l��z�es�*zG&�3��ە[�Kf��w�kN���ϻ�X�x�>�'��bj�(��E
�<s:���E��]\U=�Sx�&O�  �S�;x��Gn�U�h3m�k�9�Ċ%��Z+&��aӒ<���x�0�Mm�/��j���#~��!uW�P���%s��.���}2��vS]�r�@:8�;by�+�ojrN�5+`q{c���\��8W�u�g^�[�)YL��0�a��9�%�O@��03���:f.���!�Q�����^:�oz�Y����SW���"
�F���ߚ-.%pW�`*s�0�$���Ӏϐ�\^?�}y>�1��Ff��lHêY����i31���	5x���E��ù��Y)�=����ǀ�;a�{f��1�,�:�?�)��G���f�����yyC�{��F�.]R���R�_�a�m���Wn�'��TD������U �M�0��]`��m�F,�n+ϊ����O��|���dj�K1��g�(!zfB���yI�[��X/q梪l�����_�P^K�����{��fc���4�u^����%�Z3���(&n� F׮��H�e��;���>�AV2�w���i7�\-��L����g��^lǅ$_�����r���C7�����0P�:��:Ѳ+����ԞҧܡY��z��M�Z���xsqck���~�-���/p���E�i���5�F�'$��'�����~��Jۛ��0�=�Ğw���!MY�����gH�#�}��g�=��tY_�t�d�y�.kt6�}V�y�o�'(�,�Lřq8E9vg�J:.�:���ﾨMx�̈���{�sʌ<7��V:!���G�r�:����
�a��6/�Xv����L�;m3�}�sc,B��e3�%AǢN���vQ�L���i�����L���P�H���o�����|i�Hq�*�0B@Ez (�!��˔��N��u@1�`���K��L1l0E�r�gHe-ڊ�_z7Vxg_#W��z����O�}�\���i�����Kc��e��+��BUӖ�/cq��ܫ�\/�|��K~�¦��)ּ�"��`������q�p0h��s�8����>D1���%��N��\Duh��ޥ�SМٙ\pSxWa3����;	�1{�<P����3�������N�T�3�&l�{�����xa�ŝ��5�Lx��qCZH��[��Y�1D�"��(�K��o=gB�S-�^B��r 0����RE�����AeD�����{O���;
 ��� D.(����e��`���Ku]�y�f����KL��k�����r�g�"au�t�	N�&Z�W;�C�p�Љ��k�~��vkt"�m�_\Ds��;�/��n����UR�q��cCDn�#�s�T�6�k��OO�������HX�Eū�	#)Jb�ثu�x^��7}|�d�*Cc<�|���GY���F	�
��	U�V;C.��]�uI3I9Y>UV�yT����cf����\nR`�k6��
 ��1�4�/��@M���BO�[����G�lBux�5�P���Gt�J�>���~u}�)\1Y�1��br=J�����1�
�9��;�`���A?1��Cq�R����Q �����_H& ��L��ȝt*�-<��"��[���L�G��Xu�q�_�g�]$U�=��Hh������TzŊ,�t�E]�4A�Y�L
$��LxVbHNw��q=r|��*f7%��Y�׀Z�|	��N�jV��1�=f�,���T��<z� 8G�w]�4ܨ0�7��ʀP��ˠ§��|�z9�s��>U�`m�V�3�T~H��Хs�kJ�1ҡW_%Ѳ�֬�{�w���ԟ�#�oe�[Rj�ۧ����V����6[�7��P�
9�w��~��7�� {3+�=��9UK��-�2�����������I�!���Z�/T��ǐ�!oM�|P=�W�%<@*C��j�v?C�!���j*�R�'r�S�>)�(Y�3�k���%E�ŷu��D(T`ef:Z�b�Z;����.��ޝ������2�af�
�M@d��]���Y���c�Q*����5�0:�^[1�fh��k#UA��Mz����P9ń�T��zͱC���u@1>���*���O@�5��]3^����H����Z���.W��p���P����o�y��t�'�̎������][ �1ot|\_\�CKp�i�v��9ϟ+�A�1�CǓ�dU��ǡ~5��ޤ��������$<w+�����LO�ݦ@!���o�kp���2+���+I�U&��nD�U�W�y��Y��,�'�2�噭1*� ��SBW�jsxR��҈&�^�n� p~�W�7I�r�M�d>D~�IiƬUg����L�MVAѣ�5��	������'>�"�V��kS���/�������n�a\xD �z���o1a+��^X�h$c;���r-�:O���[{&sPvp�PjnY�J/X#%c�r��/��""���W"�a�sz��̡G��%���L��Df��ḧx�SR�\��M3I	�"�m�ǫ���Hժ3Cp�8n�;�6Z�~"{:���B�J�ڦ9Wx���Ґ�B\���e*��� ,���� чh}LƓ�-��Ǿ���Dls�����Jk�:J�`V���G7A�x%k=L�pyT�U�ڛʃ�5ʰ��H�n@�7�AϦڇoɬ��)7l�+�\+Xvv��Hw)��?���K��yvy5e��?0a�;���5<�q<6�	B�6�q���O=t9����OQO�%��˰�M�md*m-Ն�׫�Q�-x�֕y�}I�o�*�������pvi����.���@q�
)t6l��-Ӵ�Ll�h5j�w��eT!���e�`��pɫ1xwŏ�X�dB��C^�?N<� �I��F����P|2<_!����8�o�����M�4]�$�9 �UԉXiv��`�J.��/&���2KY�t�����T��si#%*�2\l�X��J͂&?���G�
 #�8���^�qj�f.[�Ř
���à����Ҝ�!.��.�P�����9a� V3�)�ԉ@�����M�!u��\[����V����T� iL��Y�&�?n��f�eB��h�b�w� 7��_�7	@�¡�\�=޻�C�ab��?,���J"濭�1l�w,d�h����ٲ�x��:�_�D� m4C:`ۊ�Q��1�/�3<���c��*�4�i��J,_��pؑ���jDp�lQ�&xݾXXS���d�Q�|��b�*X(]�40J�+f�k�<��~�iw��f��M�����
564�\\ �`��ar(�ɼ���K��/�-1!��𾅋'#��I�����!_��A������]���u���e�������:�}��y$R�*z�E�h�d�2�E��di�C6a�ش��eg�l�y;�A8��S`�S����8.���p���RҢ<���&�c�Z��w��j�>���_:�_(��R{�@J$Hb�����8���Y����p��y%#e��������	Ǉ%�����~����|����|L$KG��-���W,-���㔺��}k\��H�'��`�$E�]:�ѭ���r]�Qevݐw��臭���_�4 �As�y��Bd8qN�!0���Av�����?1U�BC��zONI;i�h�����H�R�:���p=��I^b�!�e�q�5��UZsq��C��p�1.�=�5|'>�����ԍ^7d0`ǿCu��pL�Q�)�I��㔫�M����q2����)y/JlS&?<��:��7ү�c=�@��4��b��T��f�%gk���,ɋ���0˘�e^�:PM���Вu�i1ص_��@�JT����59�:��y(�GB�ĥ��� &����҉����"}g��್��Lz��8�:�\��F���7�`!���#YΠ/%���O5��;�X�F��<�W�<)����v|Smc~�[ls���D�.��z{�֐�=��ːTÒ.s9î���`ܐ0��r�����g�����wZ-)=X�+���ߘv7����o�k^�24�٬I�R��W��n�UE�;H#�!���8��D���5}�5����B��ԟp^z.�Hg&Xu���BA��mDu�L)�ч��@����Z��]�	$�Pߌ[���\ot��3w��ש_f5�D�Qœ�e��6�� *թd�H5,�28[ ��JP��y}�	�&4~GJ��~� A貔���<��r��BO�I�_'��M3�0�|�ַ�7H!�+�7�o���%��32N��k	:�NuU3���fÂ[ƀ[4Um!�	��8�A�1�,SR4.�UE8|��O�~j�P����FA{���K���2<�����
=������\���!�K�P���G�B�����*�V�Z���1I���>��S�˂�"1��6�7��!#�!4����:��M��Gݓ
X�J��D�^(��~�#f��#��`RsR�P��y�+*W,��� M�{(iXG��FY�p~��O�HgV���N��+�/�T hƕ�m1v��C�9�E���v:	����eAބJ�Qlߠ�������x�_R�����2w����˃���g����V��ũ�$��Oý_:��_a�m�y���Y�	E�ī��,�epW,zPiQV˧9��J�;��N��u�H�a�U��Y��.�\���4�Ӄ��t�[��y��d^D��k��J�� �hQ %�� ���pu�>w����� p�)�s�aT�l��J��{dRI�?*S4Y������\����������<��q�&*X�[�d��%��Z#�;�A���ũ��'��-��jE{�p�]ߣ�(l��[Q�P��2ʝ��BN?�wə� �\~x�B���fmmP���8�c�tM�rK�Q&�E��>�{u+/��<sH�J. �m;CM�H���%D�]�K��օ�v���m�B������[�?_ط�wW���~=B �ۃ�R��ch'!#K^�'��R�'��j�U�Tٝ��
W���Q+`�hw7n5y�{��]��J&b�m$P��8�g�%�&Jۃl��)�/@ʆ�$^ĸշ�(���\�Kt�(���M.��~,���~���|z�Kk��t��u�w�@�y��h��Lh�sO�#�9��Z��`  �?T�k��	��e(�1Y�!�r� ba@GYn�כ�!��&^���2�	ZI,�����Ya:훇�v�\�&�y���� 1/xN���6�7V�z��)�ݝVz\H5�r��1�k�a��L��^#�-�o�h���^<^��<61�	&��$߻�x���2��&)�q�^^H&��]RYc�G���,�/����@wvFlٜ2j�Y�����/�<�2-D�A�.�̏�!��J/p��Ռɍ�-��EX��/�!�[��X?F�&�"�7�����lZX�^���P��Q�ԓ��M[���W/<��Ɖ᥃E���I&>��;�E�V���(&�]�$m��0�����L ���<���t[�a��-�+��&(KY��&	��  �w�7�j`Y�#���(�^���F��_���dr�n`�aهҖҞ��I�WmFN|�KZR!�B�������{��v����㕔� �Z���,��6=-�Fi�B;
��&�p�S�?�wIx�2Oah!���I��8������
�̱Oc��;1��������3Y�(�mG��h2���f]��Y��C���A�OFc�wpy�?oE,E�t!��-~N!�}�O3��?M�ț#b#(�������
���V�l�/���w�yl�ў1�if&
[|j���8��0AX���d�y�$�}�KR:7Y¶�*�if���B�)�ܘ>�GS)��,Zl�-��u���[�ǝ���7�K{D7w���2�r�ܺ�En#��#d�g��2,p,V��=���jEg��I+��-a6*;X)Q�g�9�٫����c�[�͠
;5���ũ	ډ��j�x���~$��Ď���xɞe�x��k��3ƞG�qc6=6�~M��:���u�c��0�޿H2K�c.E޷��v��a��?�B�2&��&5�m�[��:�ʦ�Uݾ�}0������Ƙ$�T�c�J�
%)���! ^a
X@�]�BF���� �hH
JQM���n���i����:2r��S�j S����&2 ����+��s�p ��[�iM��Xz�!&�l~j��ʜ=�[9J<7o����S�F�
XC넑�<������R(
�EL�2	Oܱ$Ǭ�t����c�N4Ʊz�a�+�.�H*��҄����Btodʸ��I�w܋�0�ț��;I[G�h�;Tv��~a5�gS�,�]��l��d�;�`�Q���Z��A&�!eQ�c}�*5�T_2`�wW���Ԑ�R@h��4�O�l#���9T���:<���y�:�'-�?�C�%�6pϣz�kŤԪ �����y��&D`��u�Ց�8NZ��c���h�:��4{�[����%��o�� z��r
ڜ$~k�Gx���jcAX^���5�i7�p�`������ắ0���}lಧ���ݩlF�-�����nù�a��~�С�~��Ð]���~���U&�ĕ#�����l�w�P������)yΥ�󹋯E2���f�c@���]��������F�� =�_l��y"g\A�r�)�=�PA>�s�����}:��#���I8]�.N�I��<.^�CI�ѫ�}�ȵd��L"��À����~JVgB��ޕ5�q��84�@������$���b%�9��:���ZG�Ƴ�r��P�#+X�jA�N�)yc鐽�NMjf�("��z�����K��K&5�#�/���e`I��|�(�3�Y7DA邫�ڀ�s�^
�F�FP3�㞿� 1 ?o��ǚ.Nd�sO<+�bp�6�&�r�p��W�ȍ��5h^B1zي��/��F�t��
!tj��Q�>k��5��o��	�8^L��?*/���2�@���(FO��I���w�5a �h�)7���]��n�@wyб�ֳ�V�E����քYۗ<D�!��W���ohRF��	X듛\��`��'f��܅2�hi�q� ݣ=HcT&�j���~����ǁ5b
)D�]r���k ��?�`��و�c$�x�'�-ݤ=��-|y������!��(�\݉F�Z�e�s���;x`S?�|lY�� �u�k� �n=�*[K�
�j	��Z�a��]��%��(�x�Wл)�8B�2��hF5P�d�� �jT�KaGR	�&�sB�mZ�N�OWs�#E`_�yw�;Owk�p�zN'��z�Fy����rz�2��/Oy�K�v�@Ʊ��X�ß�˞%O���2�C�;�or�#�C~�Y7p1��Ǫm!o猷����p�S�gT���?ѻ��x�F�ҵ��_3���(��n>�R���6���5rG?�F�QJ�d�[�S��%�O�FN��!aR�Y�@����8<88�tgQs ���qf�L p~��t�qj�Ո�b��44�����D��PWx���r p�ո/c��x�EC<=[7�T�	Λ��x�p<�T�o `[���:B"ԥ����u�rm��0B�8@d���Fm~�R�.?������N���K��@��~y
��#��`�'uR�F0�����h o�I�ǭ)����(��SՃ~Q��
 g�ٚ�;O��-�e?�rU}�,�[�s�@�e�D������H,���!!�����.�l��H^��B
RouMhkxs�Ў�r�V�f<��dgݚ���O���	=>�'V`�!��\\R�J�!��i?%K]�hc��5�=�s#2,��;���o��rA[��-G�:�ɉ��׆�%[ň�a%_-��4� �-$�oU80g.ZJ�TF�F��&�@�&n���n�M�Rr��ʵ�Y�S����T���QI9Z�t�
;�Ӳ�]��;�Y�Oj�x�x~�O��K1�߾��M ʈ���OX�?c ���h�r�ݶP#��.!�=� 3ӢMo���!�p#���E�z� ~�Q�N�#Hj�q��o�����^y�W��owф+��B�K��z��x��@%�_�l�*��8��,4�����m����:9��#���-* ����CQ�G���!c��@9�^(ſhF9a�� %�
/
K(QC2����/���&�1`�C��3������b��g�!�-R��|Anf��"8�:����W�0�E�;�no���_�ﰰ�}N�l�).XC�T�fk�%x����`��a����A�&�뗟���a��*�0��B��CAJ�,��?�G����j��Ǎ�ح�$(a$S�Aw�,�;S�u�Y�]&��,�xO�I����d'����'$:%?j��#5uW��C ����7� ���A�ލ8�G�f����2a��(� �^RKyW\��M>p�FG)^�< �n�W�I0����/,�.�~��D�V�x��C�ܲK�7"�΍f)�7;[��m�z��k��<U�N:�-�eO(�z��`�U����}S�qza;Oٓ ��\/Ay�d��ᩥ��w���"jY��L�|�G�N Bop�2:��u��.>�f�4{����#��_C	��j�����N��ڍ��u�dݐ��*�iq*딯�lVWy�x��H�e#���"��֬l�F�C%��O6'r����`�!���B�5��R�ry a�����s�>w�m�[T��NQ�9�X�o�'�I�@I�K���:�lb��ދ�����R>���	=ʣ�]*ECyP�8
�^�e�tD��B�68�wEp=Ğ������\�� �����ֈAEE�ߥ*��p����5vxJ��a[,����B]HYl��'8��'��
�)��WbF�k�9��Ii{����ٗ��`�-�lp��{յ<D�s�8T6�4q�3�9� *�Aӹ�\��m�5e�;li߿ĐV����4��\9��>������b�
e����ԃ�cg���19/�oY#��̿� �
���dॏp��+Z��Z�j=N�*�����t���Y3Oz�:5��i<��h'8!� l����D�{���oרҫxTq�k�Z8��E�E�R ��tT~wԤl�UK�tw�sk�����v��,`�P�@��P�mI �w�D�.���G��\�ߕJoc'�/���2�޾�TuK�D�()��Q�|\�,*�){��D$�H�hɌ��|���X��QM�Y74�'�-��L�|�w�<b���������0��iء8�g<�ȱ]l�&�`&���xE��cu�N)\k���Y�Ǟ6X�,Dh�p%�5���D��cȢ�h��;TXR�%�yBMU��M�8$M��l�^�<7�����fw���F���ҋ}(�>@W��C����{	���gy���],�(�9�7�ʱ��%~ ߈dwL��]\|䏷��j$} ��H,��6|UO�+�cc�=Y �2O�}m&��\��m��%�*?ч���N<�]i�J����VG�#�C.X۾M���.�L-H�=7rC(��`g�@ܯP X����� s&�&�龀��7����#֞_qXN�2�4�#����&C���l�=��5
��-Zu���Z���C����9���8C�ɩyL���cY�t�3"�?���#A�6��6:h�8���5H�ȳ�h�Ϭ�X����s|C��>��M���[L�dO'��<���N��FCͮ�mwc�D#��(np��r}����������X�(F�C1�N}rH�S�:X� !����5�N�˞qhx��1׳3����܉���h��0�����F@!T,J BPj�� W)�:,�zנ`Z~QPՈ!��ޣy�F��_��f����v�&|AdA��T���er~��D��V�̸�H֔�4l�T�fWU�0�x���K l��%�'P�f(��43#�T��� N�����Q����!;AI��~�RO>*�G4L(��a���F1�����膮ڷ�=p�(����S)�>w*
~�|3�ɥ���udf��~F<i@5U�:n��r\�7�,;C?��N��zlnK��ן���t+nط�f,��׍����j`$�;ʫ���o67wH��Oa�y�*��o8��%j��B�{Ԫ��J���T`j{�����K�]�x�a����	J���D���k�8pi+H���Q��S���E/ΓK:HI`����M�c���ᕢl����E��h���d�>��'���)|�9����?}�v����VYfm�W�&��a�r�.��a5�k�5f�^+���7'�&5Y��TE���O����p���W��V���Kl��P{�J;*V�[=�Jh��Wۛ6 ��hԒp�"O��3�R���k�����@�����U�ɪ�i�jz�;�k�:�w
����j�����������M�U��5�(��>�+(wR#����4j�f��I�8@8_<�?��$2��Sm�W��@���8��9Bc�rgP����Xn#�&c�����Q���ࡢ�\�@@0�%,)����#�월���+����3XZ!,���&bQ���z�,%�]|�WJ���a���E�h
�O�l�\S�+~a��&x�\��a6�
vU�mU��p��{�w��)u���wp7��U(��ѯRc�mu�\tks1l˹��5�����~S�@�zHb4��P.=�|�㷈P���+[v:V7�X����c�~�M���yR��k7%p��0���5�� d3ڙZ0z�૆�	K�_��]3�b�q����IVa����%^N]�L����Y�8�E�v��y���l��(rG��"��'�kdI��b���*�}Ei��wx�* �J ��0��J���%Ė+�>A��;u�;'`
f&�1��ӏL�n`�ϩ%mo�%��(�����r=�c3O��"Y ""�[�Rɟ~���J5�������kzeG.٤�ƺL@WO[�լb�3J�Io_E�z6�j�>\���|3V�#@jk���sv�8	RYv�ͅQR����Frb�f߉g+���^�^��(&�d���U&�������Q�7���m��f�������Һ<}0e�Gj�-B[r}��Q�G���鰷]6��C$pq��_xC��V����N�X���k���-I�����e00�|!xu�1TU����s��bI�8�Rj��3�`�f�J�j��,�hπ��I����`��k�<G�`1���t��epb
�M���Ü�h�vo��G�F�o�+rŘ��քܣR��Hp�7���#%��7���@A~�UIq]�᣿5�eU��3����j�}��M.-��ɒ{��pU@Ev0e��[�]&������\�2:�B�l��`��=�c�U
�=��g�
\�V/�?��Im��U.��uBb��
J�|�@\c�L�HG� �Wn0�A�Q���fi5p�Ez?��`)G�,���3I��l�_d���t|��ڨ��Ψ�8K6xN���h?�L#ر���	�	�Z��:^��%6�w��:-V���9��L(ΩY>F�����Zﵗ�T��������Y�4F��2f-�s��o�y��p.�����-Җ���u9!��*��	�؉��s�J��K�fTo낂'W#8{`WH]N����E10��������o�l����5x
PS=��Y�A�w��_�
;�r(����QQ��T)�{5U��Iꓠu�Wu" U�q
N[���r��Z;������g�nE���g@��]G���t*c�����fs�[��B�U?L��`Y��fV�am���s����F�+��w�����ի�s���s����Q`6w���Ή��8~!~γ|�����˿�sJ�7x��\�M�%ڧ�#ASy/��������U��"o��CX�EҺ/��O��)�:�z hm��2d���g�$M"�a�j��2�qm��O�qM�w���V��{��ۢq���	�2�?���a�-���������H�ʦ���IR�<=&��JF*#��'ק� �����Y��$6�D�2SCX�Ҽ��Q���;�č�_�4f�X�qƅ��f�5���[X�����'����^�m�n.�8lػ.łH�����3������T��v��?]�XsH��h��:�-ᇏ^�����䯞Ƿz���Ʈ�F9}��J,c ����W_!M�}���	+�H�,f��I'��TF��l��ju����]��T4�ŻGSOi���g�`J��*u��wz&�{�>&�A�	[b��W	��s�8j�=R����r�І��=�0��2Ϫ����$���&c�x���lJ��ο�֫�����8�|m���s2`�8�!؉�gC�y���'}}7c7z)�Ⴖ�	+�})�s��~��j��S�tu����/O�W$��k����ZR��k�Y�Ål�;�^=���\b:�uE% 0	�k������+����,l�u2�'�ͫ��<�-��(�&aD���gXd����wh!�o��lIr����#�`#���1���)�Xjz8��k��h�ʈS��#�RV��\u�eP6���V!�D����A�>�֠E�y�l�b�iߊb2�`�u�GbW��L�����G��d�����'�B�� "Ǯo� ��6�Q��!�Y*��G>�@3�� ��y=�◞�	7�{w���h}S��<���Z��}"��m����][/�@
�M4�ufF?�]��m�	Oh)�Bփ�oF�
��QL�C\�}��Y�6��T�c¶�~���`6u��gs���RSὙX97mǇ>���9]�2�h����(�hZ�E����D��*�RV��>a9(�j�O��+>W�|~�,��K;�ܪv�!������&Hs��2�eM]������3�_WsC�P��]��l�4�w�"�1�mn�=�Ù�Nd�Ӷ~����������ߓt{O#f�ڶ�1�!�~���9�]<�#m��n��$1�7�V�����z����siE����AUSa��[:9~�j�=�S��@�� 31C,�B����0��[y��	AZ��K�!�+�Y����֋F�a˚iH�@����}_��9>�\�$3H��|��](pڽ~�r�U��o����%�zA��9'�MBj;T�(�)���bw� ����נ�z�����לܤ���Ѹ�ps��5�q�f��q���\c"��Nl��a˙'6��^����Su0w'�i��?:ܺ�)���0�/�Y�����3՛6�Z�x���I�כ�n���~�rԇ*���@x\��uu��j/d���8Mq'�`#�����;X��>&��:���	���S�=U���W�}��tnpv��č��x�� �/ ?����'���b$<2�<˫3�N�g��}�g��(U�����,�C�b�k�&'X����^˔��I���� ��d
�𩸮�;��5xҡ 4y���|�sD)C�m�l�����K{�){�F�<T�%� o9׶�����������>�Qq'V/n�w~"0�"G79$��Oc�s8~�j�ΰ6��)Jm1?�ԕ������n<&P���.������Wj��T3�9�g ��-$�ѓi��It�����LC����D�A��y�;b�b��}͓������P-t�nǳ�F���ҚA`-u$NP��!�ŮszP���t}�ZzX�6��g(oZ�PpL/M��S�z5u�i���o(��nϭ�mҁ�|X�/�������F<�h33��4�2�(�T�1�u�'�/�N�4��yIfj���u]zD�E�C�S,��v�������*%�}V=e7�/u�j��[���[;�l�������<��T����ɘ��z2�H�q6d�`'�
�������n���k>���G�D��-��E�2��I���_N* �.Gs�S�,"��Eµ'� �,u�o��K`�ָȽ�MQB:Ʊx�62j,��k��AjG��Gz!��9I:����A�����\�	#�zu�Ij6J�u,m�ˇ��&'�v��wG��>�ˋ����� S�@���Ƭ���~Y���%��W48ݬ+'�9bw�O����v�H��P���J?�x��m�뽂�6__H%�����5M��h����-��`���kMzV;`��~�O�5!jk)�"�^�Iv��j**Z��&s��m���?C৓��Bs9�Rx5���Q�8U0��~|�����XqY�룃C�����B��"ǹ�� �����,E]�%2��&l��#=YG��ZX)	%a0?hT�,s�~�����׽2?>1��Ǎ9�Ւʖ��)g�4�;���_����*���3��Gd;2ĳB&Vz��
Gb:��s�"ߦeo$�e���Ŋi�sF����w����ũ������d��Hr=������'��H�+>�νz��"��y�,cy�����.��	�Ӥ�P���zVA�6����q�>2���$�v&/?Kh���)�kD[ �ʷ�\��Ğ��'>m'��d�Yq�a*�s0������J�R7�����N �iT;�_�z.(��__'�,�FP>׫��rb�]较���b/2�CNjY������e�r��h��@�E���1�#H�0֧R�G%�*�Ƈ�DCǚ�6[�g�`l��tO5�K�s�m�Gc)x|�\�(ք�Vl��"<�G���ԛi
*�[�R&\�]Ѻ׫8��'���*'� t��r�e=��j���1�z^,Yi7Ӳ��+o8J}�(��p@(/>$Vpi��Dz��l��c���W`�f�؂��i�6�&R�k��p}�[ik�g�!��m~!a�_]������3���,3�(Ph��B<��K����kx\Bn���������w!���n���u7Uŕ���=- ���6�*!�X�]E۵��x4{7gY�̭ȿP�y�-��.��˲����22)񵷭�.�9�(�{ :��zFO���|ES�=��42�/��n��7��)O�V���:#��sm��
���7�Lu�;>��E���M��v���sNPt�����/Dd�������`r�I_�Ugo�$�Y��ا6�>"k6�3���;��?�q�Gxuv���U��R^ɽ�^�Q �8/1y�+�������W��@_��c��J�{6~����O���e.�S|���xG͐O5g~[ʟĨ��Ơa\g�.�?'�=���ao$��6~UD����TL�%����+�F�pO7�e�eEY$�8�=6��X�_d���SL���E�I^q�z�1�iI�C	��ތ9�0�B���s� '���R�JV] �f����p��CD�ML ����U�8��& �7!�$�*&�a|�/\����ֹ�/[9H��Q��s��?/�V-zg�֯ӣ���q��R�p������_����KC|�m����-2��tU�>׷�q E���mS���+:RJ�2��9��l6Y@��P�G��`�V,s�}�U��@BJ"��b��?h:5�w���TG� 9o=k�����թhdS4�gQ�I�V��o��=^�l�"�bq/1�8���#�z���*6��M��0����B�b�.�pcDmK�Ct��.9
Y��i�̷~%<�-(�g���,��<���������l3��8��[���إޗ�n�7��>�}o�:DE�6K�j�\�*���!C�3Y�,!w>o-�?�3 ��p�[�(�{s1� 3c�[�J�'J�#�����o��Y������G�8 __Vc����d�*�I\��V����L+�+�~9r���-��è�<?cAh��beU�B=�@�b��]��&,!X�%����i��(��ݥ���Sa��Д�O��v�PB�cI�p��_�>�h�T��<�*�Un6`��G���:���"����U~���/<'�j��y��h%�����מ㴍�Z�"�����c��=��ڠbM�<k���$21����z���?|��־̦"������y��g-��?$�؜*K�5ͩA��E���C�Y_IB�����'��`�dR'<<м׼�~��}��F�m��s�zf����搐��j�k�O���5�ʥL�,�V����68z�Ks�Ƃ�[.F) "|��۶�����oݧ���b�ueP/{�p��]�u���RvN��=F��C',+6H��>J�^�qvŽ&���O�3]h��x���sp;dW�K-{.kr�\�v-�N1P��wȟ�]��P�wC"�d���#EJ*�&׺��w��P	�6��a����ʜL	�5�JݚI��~,��<�&�X_���A�,v#�լ�<����R���?�p=���8jAw'u�V߮S�{D�YB�?-W5sK��5�]�ؼ�	�ڶ&��!����?����;�v��f��`:�BPGZ�@���z�'b�n²�ɒ���Fδ"�;�,Z@p%
K��/��a���h�;q�)�O�!Edz��8Ō�b.%�ũ~*FV֮k`#K;g[<�S8qMB\��6R��;M���J/��B�6�ՊV���zB�⛌`+�����n���iWm	Z#�R{��湔{��VQ��Z��C�R�=��U��#��)o$yz��P�^�L��Xir	c��y7����0rCVI�WQr5�u{��K�>&]a#j'�aم �/�۔|4���u`R�p`YѲ�xz��� �S=��OLF���I?�2��x�|P3Ҫ?�g�&�I��B0�=����bTׁP/{�heBD�#8���&#i��5gV��'=�T����a�b��u�7Ď����^6��;ыd��."ɓE�;�m�#v�2O�e��S��K�6���s��D�w�[-��|����d&�r�k��O�J��L,���x�0Ե���s�~O��Ng����� ־��fء��(٪k)��Q���(���{��W����"o����5��k� Т�X{i�}��b����`d��eu�q&)�h��Գ��r T��.�����Ǣ	 ��Y&	�'�JT���
�o3�g���A��2��CȾA��!FSS��Vɴ�:���C��vw*��]���ѹ���Ex�fmU���*�9A�u	&�Q�J Lq�h�Gw�M����	��xݴ�ʖ�����f�ѥRqC�YԮT�f=��σ�lg���c�ͰS���@�G1���|ϥ�-������b��D�o���.4�r�Z�x?���G�հ���a}j��T�����5���D��t}��'�{0dH�iV�ƶ��t�C�)�p�&ɤ#�,"7���*�"$����^[U�������;m�<#e;�S��]7�lJU@᳦�|��KϹ	5:��Op�cuC�SF��Ƈ�p�r:�m|W�y #��WW�"��F�l��԰Ѝ�wO�z�H���@+����\ȱO;�����x����$v��yd�k�a9��d��vxgx����K�\�"�������	q�n�r2�4��w���W������tm*.(�$ӵ����^�I�.A�4t�О�L*P�u}	�l��Zp�� �f%*�!c�b�A�?�$���%��������gp�)��َ�޹������孥�P�#�r9���R����?�ܞT�Kcd�n�Ԯ�i��M�_ED�i��L�L&��~i˖�!J�d�b�[�SM�/��-ӫ=�{}-5k>{)<�U1�8m]#��[��Zy8�����d�� r�FC�X�/v���m��s��,�C�u�$����]��_AO׽�NSd�:ʬ��Z���;�Nj?T���� f9pZ-�n�g��!P�ޛ��� E�0g8>Z�]H�t�At��0���B-����{�'��L�^�<Q��T£�vtBfu����*g2���~s���3���/��"D��N�H,��ӔL[��p=�2+��/lPf���Q#�5Nm��2�Ӄ��*g^�R Rj�{^]�΄Y�##�w�N|i��>���AQU�M,΁
�Hx'R���p!�_��=Ė�:�o��x%#Gg�܂��mcFj�F	�Qˌ{�9UҢ�n)�o2>-����ռ��P�"e���%U�sv�]�X�-:W��5������M0[�)gQ�$�綢��?��TV�H�N)�`�jX����:��6L's�k����*_L��A>3c��Óz��}��pf/l�c����ʷ��m4 ��1^J�R���n�+~�	������&I���t#�2�F��@n��H�f��"1=�;��d}Cm$�k��˗��$�s+�8�!�r<FY*�=ɦj���$<�e��U��Nc�8u�,�\獤�����"�N���#�B�;]~5e���)(iЭSG�s����s���_4)O�_ï|��$�J���J�TΒ�N�1q%�-��m�M�$-Q`p5�W���4�uYG'��6�u�� ��6��=\~{��:�p-)cG�����X��Z|�O<ה)��ϟf[�n9��=܌ ��f�ƾ��f��K�KS⸺��A�6���=t�~�'f���r��x��Ke�Ж\��5	ˊ��8`Vt�4��|���S`���1��w�.�4~s�{�4F}�0�/��_]�h���1$R~��W�T���;*A<}��� E��#�ns�%�����읚_\���ۡ&�S��q=$L-��7��H�6��󥵃J��ƥ�7y���t�Z�-����ۧ�-���N}����۶�>�݊��F��G��ג3�tT�̿��,�k��PuQu�1ث����#5Q��ޱ����P�kE�w��Z]�m�*�_��O���"B�.�|Hhi;�C�r��D͸�7�eS�"��#�ߏ{ճ��48�ĕ�S_��-:��^�y�	�)���b�ڶr���LQ.$3�=�y��
��x��L�1��I�r�u��u9���(��I�=�iq!MvK��Ff?�}�嘙���2���0�Y�����$��	5��T���A=u�Q�}_�����&�_�`��wk/{�82��X�k`1�*(���1�/��eB�c6A���fQfSL��||��;�{�ۤ�˶2G �-~���:�^z�@M(6>���F��S�PniPJ(bwy;���4ҷ�1m��F%�9���R9�܋�k���M��iO�D�U�c��U[�FI;��D��N�%yG�7��C&�C4N�Q��tZi)qY��A�:���N��i{zP����u�ؒ5h@��C{��%��������e�1n&�S@�
��+�P䱯w�
�������n��* [��@�-�ad���� �%(;d��N`irB@(1�	��������l���O�f����}�0�x��;�$�\ɃeR�n�(�#BS���+։Y�+�����?����_19���&S�{a���35���+I��ܻ��S��}�}�+[y4R�]�'�����xz�rׂ�}���\5\�s�`�>��#.�$^�C� �LpAܿB�}��d#1J�p2	X�c�U@d�� ^ךB]� ���N���$}����S��*�������G���h�h������	�.dv��gN@����>�l�F�o��w�W����;�'��9�ԉ?o�|mC��5ys,B^�¹�(�8��(W�
���^��5����0-PXcJ�?���uI'ho&T@����Q�q�H/�F#}�������M9.Fk��9{]%���vj��?6���{x:H]��y��CoThݳ��-���I�[��SX��m���$�8�e�:��O�����T#������،�ܠ��� �0����6�h%N�-�GSX�&�	�Jz�:-Nz�*���K0��`c%/������=|)���U��!N[�5[���My.����Xx8a)Z�����o�<�*Y���oo�z�诗��Z��k��MM��
Az�gE�T<�G�B�#q&+O|���t��%8�N)^.�`g�����&���>�)CKp��:��E�~��&J8�NO�HbB���cqq�șx��@����-`il�Anx`�û-i� ��b�T]귟,�D�$~�
�rl��N
�Z�7�ܸm姦ɐ�;vD��k�E�e��.��2n	��e�j�;4�r8�ގ
Sy�D�яE�Ok)@�[�k�E�SY)�w�D�Jq���z-8D��G���B�J	���/�Li�豧վ�@N��7O�6��W��,5�k4�����H�G��.sQ�J@�fv-���6Wubj/j���qX�x��y�&k2K�3(�}j��<���,�}��ii�Ћ�^�f����țz���4�#���4z2R�)�
U��יj�h*6�}�v�A�XA���O�W\��5�FD8pG��/+*��iE_��."@ICT5M��+KHݦNTÊm�U���u�����Փ�g)���>b��O����p{�x�?y��A�u�SҀ�8zF�`Օ� }u�O=�m�E?���^�Ef�z>,�X5`��&Ѝ�_�Vk�	#o�,(E��z3���Tu�Y�1DNWϢ������o!po�?��\�"�f\�����d�%)��	@�D_)i��T�MJ;ޝ"D��ة�% *�Ԑ�ׯ[/�˫��ZH�P�����>��FT���	@��RN��V�<kw����>�?4tx�����]�գ�"�|�?�Ѿ(���{�:$��=z�9���bq?�U|���Zc����+rO6S���2�WM�3B����IT�Gw�,lʟ�p�V�e���A����E���z�Q��w�%,����4�
��a�=Z��-K������I�'UVb�2K�P��X�ϟ�30��$�}���y�6��V�@������?��)鋏��^�8�q���N������H, �+R!�Y�kE�p
����I��4�둝��@j+n1A&��~ �03Ck�<2
�/xoƵ�+��?%���İ�]{����}P
������e�,�=��� Ʈ�����'���f��] ��:@M�#�£��T"zP��g|')y���o�\7*��i���N%A~*��S�\H�4�+�15��C���O}?�\ͽ��n�au�?1X7i�BW��*=.��p�ޟV%6z���^�@��"ܦ�e�X���ƍQAӺ����I��"�Cj���C�ܨ�F�Ӄ�}3�@����L��W�$V�E�C�A/ǀ���N�æ��Yf4�4g(t�������G���$����_��ԍ?)�����U�����'p~�N�J�D(�DK��/i%B3;�G�s��-+!|��a�M*����}����Tm�U�85m�r�����|�}�~5'�}@k��n@9\��
$�Ul��b`�z姥zl��!,�>M�S���:~XT�ɛk[�%�8_�K���)�0�z�&lL6����h��]':��m=K)A�-�n���OM�ޭK_�P��������7II�<RL�V�ܤ����6$�Mq�^�=��Fқ��l{Y�gֻ�X�Z�K5r[\� I�E!�90���^���l����3ϵ��@X8�j[��I�XA>Z�4��ʠ����m#�7�,Ы[A����ν�5�*�8�3[���ȗ�j]�υ��	�u(-�o�rv�q���w;�SrY��R�͑�Vgp#!���,��6	(��!.����-(ޠ��e�Y�CX��,����$N�y� X�J�faZa:�^��r�r�#޶O�>�j�}|�Z�'ȱ�[z�>�B��ST�w���ARM���IB����*X���N��lo3n��Њ���'v2�^f��ɮ=����ޢ_ �+�l��iիh�B@yP�OIׅ�����)�y&�Z���;c
���ϲ���Ⱦ�~���x��u���S?��M�f�L<�ѿ�Mj��I�+ڶ��o�Ɇ����O������7��yC������Z1nS��g�
��Y����t�o�6QH�5�_�lY\u�/�~��	*�/�q'�m.:G]Gz6�"{�@3�S�-��;<���o:��1���%Ƈq���!Y|�'�9���1�_�A�IEUjo-��2�s<���ڑ�H�B3<n��Na!9��gsQ0vg���^z9��a]��fc�c
���I�$)2Y��]9�Ri�r�[�Af��4~�)��L���$��G��k�]!w��	j�n�۰�.���u �N\��y��QPI]-#�υA�ܩS��.C��ގ�y�nZ�S�4.Zz� �V��a:���~d6�gj�Z�i�sT�UM=�%5qn8�b��J{����^��$N�����j���7rl���w�$4Z��F��c#@�3�t}ci��z]�ʵ�F.�\r��M������2'�39�|1j�Aȋ%���|��V�P�D}D����?��TN��8<|q����p�OKY�w���
��"�Lv�{��xc0�BXn��ۇ�]?���Bvk����_�#����L3ݵ7�u��I���`� ~�<S�.L�:<ORȦ0��1;��v��_k���`�B�j���T%�������g��ĩGz�_�o;O8H�ݯ��+fW_FP,�OSQj�W�f����y���n��|��1j��z���T%����z� ht�J���Q�|�6���`���h��ņB�I���STW�XkJ��{�mwuQk�țڤ ?���W7n���Ys�����%[���E�&cG�C/j�î�*ō���X��"ʕ.?T��!R�@��y��w={��֫w.w�2�7�	`��R���	��#�+r��!ۆ#�`*���8��@�b�/��,��gn�}�7��.�) V&vF�R#T��	����v����<U�Ǵɯ��h�_q��g��)��3:oU!�^o��V�1ѥW2<��F��u���v��ȧ�8�8�x�����dx7 �d���2���d����� %5��˛(���?�{�i	�!������u��ݬ8!��a��oYW�[�yft�4UHL�������NE��R�eӍ�w1�#¨p�x#��\�'��&��t��ѩ}us�\�0�p�PG�T&�p�u��7�?Q�q��e�	�>F&1�@L�j�- z�#�G�
�0��X�q$k�g8��fC���$��T�W���Wѽ���L�����di�m� ��-P[����s��h����T�xK��`�V����S3�ojvI�Lr3XP���Y~=K~�v�rC
{�����׮���͓���0Gh�q��8,f�2��`�8E*�{�d���葥�����	�{�UE��}ű��L�{��)�Y�h��-��<�A:�p|�Q�V����^ʟ
\J����^��T+��ʘ�
Ёfz� �����!0Y��b��/�=̈򁊃�-R�Q9*��G=�����RD���`�@(��^�
��������4���W� /(U�Uك���4�o�5r���G�	�/���F�cb�����i +۱��wֹx�������j5��>�0��iΦ���v�{&��_��	�v�%�FU]e:	�԰��>?�h�@�\a�@@q3,�Jf�PR�z|~���E+3�!�q=�?5�I`��p���a�\��q[���!��פ�^ɒh)%a�Dś�Q-c�dy2ʻuN�AL.Z�
��٫3b�L�e,@h��e����:�M[3�;���MKR���63$	n����טD���C������Ei�i� ]ҁ4�mm(L������ϓ�%p�e8KLll� �H�����m����{|q���+��1#n12G�;d4���Z��GN3M`��V����ÖR��Z+���w���`��[đ��0^m�"?<6p<�V�g|�%��*?p�D�?����W�\�%�`-��Қ�E�@�0���jL�P�N��;9���V�}@h�����$�o� T�=T��H
R���\�$q��'�.���}g&���S�%k�ߒц�q:9û%���L>C���.�:�.�V^�dv+�%�R�f�O�Z�K����&UY,�-,���!_�s\�[w���=�����V@1�C��W��h�U�?R�E�Ay�3�w��ȳ�΍o��r�x���=X�Ҳ�׿q�8�E��.ާ�	�>�!��
����n���F;��V	xr���L������/i�!:���O8��#��#\��BJZ_��a�
�2RM9:�e)7Jj��l!J��$�+��AS��w�}�-��Tk�k{m-ݶ���v�$v�d������<F���[�4�mS�r�C�f��K��/�WXڹ�b��!���ye7�~�;|�W!H�R���ӯ*���e`q��,-�p����XY2j�	�q��NJ��ଃ�O�%QQ��[� �`u(�=�2�#��Sg���+73t�C�T
��w������%n�'���q`&N��í�|T
A�|]h**;��;s�����u�jnk[X?��jӭ3ж��k���[���{�0�5V�?���SX����|Dٳؠ��I]��df9	��Ԥ5�ˀ.��*�:�s?o��䃘�,���f	8��@\�?��A��W��j='���餛XQ�_Z��-\�l�P&9]��"�-Zhsǅl
,m��櫹�S#�%�W�N6s`E��'�"9H�ڟ�)D��q��b��3;mS��	8z�����m��K����8ˍ4`�VM��26 3uD�gk�k	Or��_�f�0l�mG�$�m�CY/��K#b��K��M'�=�Y-!�������m��� #K�c������j��f�U����-�#xV4zh2����`x�X�o��a��hJ���Cb�ai�\Ƿue�b��{Ea� �U���|:�5�"�HbpL?�i�IE����Z�	Gi�!!{D�]�d9>̇z����$P�!dyy�ݴ2�>���9�"1Ľ��u�)�k�� Eh��c�g3���pqXauS�u5���e�֚e�Gd�Sy�. 
��5X<��
\����%:�G-��[ٙ]d"�,�Ìs�焸G�b�|����bjXK����\F�Y��LI��7N�D���X��_$&K�r���ېXz�¹���P��"q-w���/w����o�j�)OX*�3�i���]�� �_����7�Ŋw�Q�Yٷ���/Z���q=7#,����6�8�X!"X�y�ѡ���F�BƁC�n�1lf@꼌�$;Ϡ��$�Oaܰ��V�݇�̫[��ВZǢ��v?���L���Z��-�R�J~f���~9�r��V�:ˢߝ��Rg��2�bC�zO6,��������Ӻ�\ա�,v�Û��w��+�^L�*�'(N�K���qYV�D��x��Ό:?�
ǚ`�=�jF� a9�N��xԇ�6�w��la���Pv5-�r��(�Oؗ�bp�3�����(��/�T��U��֙�A���1��Y�
.��q��άwθ�B���73^(݁r�����?	��g�f�/�LH0%�&���D��o!/�&�����29�וa�Q�3�@���pg���H�m�ε�=r'�͐����&L�#�(�5f �T�� d�7&��V"�S�<Yp�^㏈��d�]�,�Y�dc;Eb�v�|A�RTN�I�w�J���Z�f�$��yp��jj�&&E[���s1�7�E'��3��:M�����[ٻ$K�����ZE��G�e��L����ۧt�`6@bdS���℃���5������c�5�/�"*��8O�X����+P7$;�EM�����/�b�ܥBL����R/ʭ��'~�Z���u6�.�\k�_�J�o���0e��ɱ��*���C��Y?�=F]�%�RO����bxZ**�W"���W]�����t�Bxq?5��úo��g1>)=���жT�D8e ������i�ׅE^is�c�}$T��i��'��4ɲD%|�
.��; b;���/c#XφK�#amdy�-65����,	{��YNy��}.R�ɋ踆k!���#�g�(��۷�y�g@�I�e0k� ҈&�HQ1�������Zٟ�R+�K=���X��Hץg௺&И�LV�W@c��-_�Q6��\Q��R����~��,�e�8��B\��G}�m�ν('48%j��x[:�߫ڽD~]���h9��lv�~����� l]���̷� m-�3H�/��mA���,l��6��K��q�P�lI5y4#��(}���%�&��B� ��dw�������ChZ!P)x�`Qψ��\0���a�L0S-_��	��xz�Z���q*��#�P��\�r֬9{�l�����2�����:�H�]/%�E��K��r�(��9�;[�9Zb	_E���C���S;g8-s��\��ՍInG��Oϫ�봬|���P׈p� �p�[.F�ii�� ���%}�d�ZUh�w*����M�ï$���>M|��iK6�
z��a�������'�M���C�<'��˿w8+,������NCMUw�3}k��I��ܪZ�i��9�� Q7��>%%���`��~A1���0ش�#}x#�<MߕO���q�߇�� �~��'9�{+(
�P�u�ef>t6���>CoFZg��ڇw7l���z��N��;�%_/؉��2����`8��i��F�P�b6�]�5�wG�����qg��*a��Ѓ��Z0c��:5*<F��˹��@��Ж��g糾�zZ̩)��	�3�Vu&x�1z8A���D�&|e����N�x'�d)\��Y�@�B���
 �+��nCt�zv�N:d��#Z-����̏e�%���E>��#W�\�l�)a�����(Ƒc��qE��'�I���wM���.�SB2O��P`�u m�Ĭ�"�ř/=�=�����d��$����z#F@e)V�~m|LRN��u����ξ1w�W����:�Uy�bD��O ��}�4��LZ�A�߰�L�4y���k����м��bi��(ЅB����`u�(`��r�W��b'YX�q����kj+!���W��?�7�ʇ�N�s>8�s�z�zfLF��$��7]'���!5�;p��r(�΋7��[�ǥ�bJp�������@_�W���}�r�����q�DS*O����$5'F�F"f��B�C�GRo�JH_�
������w�JBA�e�?!)H�hI�Nz��1m��O���,�H�E���fuQ�W�]Rf�sE��jȦ8԰=�l�WLK��A���t?�q�*�1��	f�DFPo�v�P�[��>7�O}w��e�0�Di��������U�ř���0�n=v��6d�&������X��u�YH�����E-��EZ�xP�c�xI�	Dt�.u�L\��1\z�����)z����63�F�I1�beý*��D��)�P5o��r�yy�t��B�*�VW��NR:������pV5x�b��<�k�`�,W\���1�B�c0O�#D3�)6֍)@�\�9�))'J�����.Uؙ��~(�?�YN��NX��TW���7ji�i�U|���K�8�#䉵���vk�w��❇��!�`챯6ų�5LW��AJ�Ne&�jdg]4���M���>���z�o�(Tp����9r��\�oe=�F�#ĉ��.n�=Q��RXq���u _���i�>9�/��.��¶40�1��M�-��W��N�o.�Q@q�`��u�� W^�z�(���f¾��l�`��$��4�d�*����n�������b]��+�9���L�؂�N��Y<W�{�;��V6K�m3�����M��ː��'�����^l�A��w�L)�%��gQ�jI�y�����8.e�P�%���zHyQ� ���w-�����4ܩ�m��������/7eZ7�7�EɅcu �WK�=ʞM:��x���㿠�7��B�++4�۪�n��	 �UU�?�vحX��r9���r�W�i�̶�3��4��*��~�RCqF����&-
�Ō�����$8��V�I	RZ#8\���N��5���_C�)��*W�7j��bP~� �p:&jN�sȒ��&�Ll���x�a�{:�pޓ*�-�<R�	��l6����s���/�K
�cT
���9._��k��\�Z'U'
C�<����3��v���T�Fo�B�v?��hz���i$�^]�D~����7m|������ʒ�$�{0	�r^�����1�}���)��m��tFj�n�a,���������ɹ���+��/�*�x�J]��M0E,�Ŵͧ+~��o#���A�	R�&N�-K�eO$�y)� �%sWdL��4���*��&�;���p|���3' �֜0�)�j֒[[�w��&���zn b�IO��]��(���C�$��E���o/��l?�O��F���0�ڡ�?���gpB��K�h*���T}�j4m������F(�a�a�u��"*� �DLR��_��/}�/���W������)�f���q��[aS����S�.�]���'�b�H4f�^�iY�aK[��E��<�û���݀ܣ��3�T�A�m�p�iG�+,d2� V����m\]�E'���~�r�U��nX������Tl�6��FP�V�y�#3�n���*��B�LFKw.�,*8z H+���M�Z_T۬���T�mB~�����k��>T�?Z��TL��Z9/r��j ��#�yB���q+��V�˙�.
>_37���˃c����f��݁��G��z<��S�ȓD����	���%���w%���.����͈�Yx��EI%XӐ����n����t$�(Ex���93�øo0��_D��I�.g��9`�Z�?���=/���⫆>� ��5��N8�%�:��N�pH�i�[�����7EE�XMn!�A�Qµ�Cޗ�L��C��� �`ӌO:�����p\`Z����̈́��O�5�̑W8�9$=��ҝ���S�Pu��^Q�+$M�A�O�Oy+`�=aV�x�kuPc���%���d��S9�Z�=�-j$W#M�h��K�����'�>~UgU|{D9�?�GV�H?����E;�U(��۩��*��I���i4d'���c�9��(��cL�	��ь���E��*&yjP��}I`[��K�I��XI���U�/R�)ч\�yG:`퟇��,�_K��FUx%�VIԻ���%=��e6�hm��1�a�,m��{�Ϯq;=�=��f�0��%�A}����U�R�=�.G#�r|.Ur>ޥ�w��/y��Ԟ���RXޝ7�
�n�� {��]Eu�XF�+�#)#�=���:}>~���0�i�kE�H#�;�3������}��P��fB�=�Z��hǰ{fk01��.��sZ3@�5��� ��X��l�z���@q���3k�*U�>�]ރ�4�#�:V<�ު���导@c�ᬀ��@�������ڡ4m]�|yrrE¶D�|k�_�8������)�݉�W#��j�����
p�o��KZ�v�cL��D��<8a�7D�At���S+�l����dzy��O�V��38ش}!Uw%���I�x`w\��c���B|=ᙬ�3�_��Ơ" x�DP�N�MW��; ,�uB��9��� ̯"��uW`�e��}��S~��5Ӭ�����5"����_"�3ḅ��G��-�P�_�?`���#���+��%V<p	u��D��|ϕ>��D�ۂy�<p���Cފ�0��a�3B���_�|#9��/�glŽ?cc¹��?�sq�l7b�XԐ�}�zQ����Ɵ�84��3JIc���Y�dD�W+n���a���&�z}2��w&���؉���nH�N�L �S��,�����[I���W|��N�������hY9q�>5���/��|�\�.^u�]���Ґl/z���PEע��-�� ���@�X�o{5�NS!d`���N�n9pK?I�j�����E� ���N�(7�t{v?���W�7�$����;^Ss 	7އt���D �6kx:s�k䂞ˊ���m@l�	0,��m�ܴ�vR9�K�����^�"�>�A6#�/b=�S��	Ŭ;d�������� h�I]=�}����b���L�<ʻ��'k߃�=ǔ��o�5�F�"B���U� �J���,#3�+fTv�V�Gw�ʷW��F�����'r]�V�'��sI㵾�)�e2s�f-�qz0{�������۟F���aH 3\S8�(��u�$�l��,���v6ֶ��e%�7hHH�v��*��˼ZpCp�E�e���
W�Z��qܨ��W�Z�ݲK���"�^�ד�k��6@�Ή�m
T$�p��f�W���������}|����FeN�;��Xwj�5/%һ�����;���ʚ�f�d���]{W��x���k���Eц�$[i]nvODK��|��
:���w��ȃ��lQ�0��������#Is��Pm�9]a��P՛=7�@�Q�o�Z�I������Jq�Jv��q��nb�k|~��nތ���ʤ�!�#E��<*#Yl���<��"O,�~;-��P�
)�����[C�h��4G*�ߔL( ��<������"����y���'�`��ui�o +�V�#��*SW@	���֟�����pK��a�����Xu�O�I��S����u���u?�2┑G���Z �������ٻ�tf��ZO��x�Op�EA{=/K��TM�������WY��v%��O�˧����u��5"]F�p�ۍ��wN�UL*y+���o
�{�N&c�.�~o���}��[c�J�g�|)�=�hCw�2��=OVժ��K$oܥ����HFĔ�&�WA�V!n��S�$ʇl��*���Z)i_�7�2#?)?1�¡��(:��a|�R�{�$DH��/�c�u<��g1M�h�е%�]�W����~�a�ψ���MP�K�~m�a�P�S��;���N�f˖>���!���%Ǉ�s��_��7AI��~��
IB��<��������I��A>�A����:�
�9�H�f)׻HL-��H �a�B�^���}�"˘� %2��Ɵ�'١���6��6��L�0 {[Ң��A�MPk�ۊ���:�4!oW��y(L�Iꐙ�6	˒Ɩ͌sC0\)�Q��جs�ՈEU��gY�.�].=�a
���m�}�f�&c�`jH%���l��s1uu�l��ȇ:9����Ҥb �N������O��l,�<�Lg��U�>W��'�2�E$+��8��>� �~tO>�o�vρ9�hK��ġ��V7����A�V�m��`(�&=���{�u��X���$��@�<�$�4L�=�[���~��I��F� }P͈W�AͥX�. �tN�du��M$�_V+|: L��r��t�"�|u�$�/@�M�E	<�g����p�9i(m�%�bW�UC����j/�Bte�5T��b�b/��j�K���e��u���~�)�:�,�}^ޚ�`�� ɴ�H8�6vh0�3������<q�>c^j��
n�J�H�<EC.��`��!#x��6���G�[��=�!@�@�8��C���es��(!�xZ�җB������� �?��ٮ	�\�a(\V��Gy5���[Y'k���u�555�H���:�
�;�����ZK�`��Ί��%��k-O�۴��U�NNi��7���K�ǜJ�H�3-�YMaϣj�����6�]��:���^ܬ݂���V�Z;F���6]�}��Ėݑn�r1�i�zo�߼6g�v�*>���,�{C?v\l@/��_,�J�Y��a����`u��׎��қ����j3��g��ݎsT#oES5
��q�T���ɹ#�*7���h��w�Y��t��t6�]��V���ӳ-�K:q>bI[y����Ed9��1�[E��d$**o�o�O��_�f�	���wOs!$h�
�����:!�,L	9��R��<�ɺMd}��\cu���6Z�7��O,�~�����f�]C�!!�t \���K��PA��!d�Vj�I��O��.��'GO�C�w���{!U�`�i�9%a�LFH<f�8+�z�G)�0>�<�b���!�!� zS&�Z�5Y�k}�0�IӍ�I�g��Dp��v��mn���Q��;?ӽ����l֣_m�]�f�JE`ƚѸ���3u}��G�uݿ��E.|�t�Tߑ�m����y"&݂Җ�t'���R;ea��B:2�v�0WE�れ�z�s<��4iz0�E�Du�C��X-q/�T�}l+��3G��-!pi$ �N��!�p)�z��X۫9>!��6���):�lo�Teۈ�N3�w�(ZY��K�+e�k\�<��" d�Uf������5w2� 94
�=��Y�d���g`����zKLö��ha�%��X�.���=� ��}�G���Kw�3�ڸvb����>�6p��	_hO5�0���c�'�G�.�"��������z������z��,�`5b[L���hܖf�2���o��t!��MV('��KZY|X���í��V_���0eC�Z��1�ٸq���-�hO��r��n'U(
��Җ}�x@�g����=Z['�Bk�D��ْ+��eP����>��ۮ�,���f�7ʘ@�~����{�3�f��s�e����!<y�;���r��y������oFjy���ULA�98��a��z�����{sϕqK`���6��=א��pY�����st����N�"Q�축��#&*=�!��J
qa�+{�_�CFzZ,Yu�~�q��J���yQ��9����{rEk�﯎ܔ�߾K=���.�l��1�Љ)�Y�&<V]�0�m4�q�;�"�<�bg
�هE3/��Q�'Ru����B,-k�v�SC	�� a�=k��8����,%��ic��[8"�Ey�$o����v���L��r� sY�61�fݹ5P5�.��N��bڎ,�O?柧����)�Db��
�a�<��5�⭅*'�q�g_�1���b�+��?52���ߜ)!28�e��u�|g�o������{.&�L_$|���;Ka j2�G�ޗ��@V8!�.�<e�v���P:�OX��:��4��Ю������-#�|��9-�|Ֆ���Ͼ�bZ����A�T���M��t�<Vj��Z8�\TT/��g]�A���<y*������u�E !S���q�����B?=/���:��S1����MCG��}J�b1���Gu��W��o�Z,���3��`pȩꆵ���v�?U�|M�o�ɡ"QZ(^u⨈���{_!�?��f�'�G���.o�����k �����0����r�l��q��F�H@c�M�M�O�) 3)�9�s����S�}���ç&y��S���"-����-UMU{3�"��,Q�q����j�20C�>B�Y� ��(c~7�
�1�k<%ٝ�x�U�M_�x��͍?��1�r�[����"m+����|�nW�=���[������Z�H5�*���UZY�p={��K�`o���#�s�U�$�dP;SK69�y��h��4�ۉBP)�6�YkF��eW�����q�Wa�2��M;�c ��p��_1T�7ڛ���^?�8�Yyz�X�=�enj�����f��3���=m������d�4-�[/VK�����.�}`q*�16���6kH��zA|	�SE9^�!�,�e��wb�=�DC"�����F��?U�c
�e�L��1��f�8�ϋ*uaM�*am[1�p�*P��	jJĎ��.'z|oC�]�p\^+�M��,�pe��soE����F%Qi�)�{nG��x�����8�?n6�?���/C��@�O�'VJ!�l�h����q~�g����zɃ�Z_}\C�X	f����0���X�P��~���
�OZk��b�$����?Q;��	xipCU�N��2h�D��oB?9Z|�_��\���l|Xw��u�Ģ���S2.[n�&�s�]]�it
�\4���4�1hϼa�_s�uYr���|Ѕ�ְںm�xQ��r��$Z۶�!;�����4d�=
�l���[7O�+f��>�4ϕ�BU֖�v�G���g���ՌK��ąC�,�'h���q�"�<����7
�4~�{6�f��{�� �K��:�P���QKBь��Q,� ��K }�Z��%J�.�[����Dx��E?/���:ˍ%(��2�)BZײ�F�;S&��%}}�qV{�j�<��W�B��<X6�S�0��6�ڜ����f\f��a��H`5�Ti[��X�����N�i�)����H�M�಩��&�8�44À�x���x��]�4�+�Vòď��9�M!�pP�Ӫ>�/-�E�����e˄!����K(��8BȃN�5?$)x��H�� ۡ���{X��l��Ȇ�)p���.s�Q�H�m�#D2\l�ْh�ٕ���&ŗTؐȠ�<������{�>�*s��� �M ~>NaO��n���/K���A�֘�8,��5�<t弮Hj7�F���:��ތ*p�Җ;����`���J�:���Mb��*\S�&k���+=�\g�{Z��y`��]}����o�:=<;�Km6�<i�\X�Z9Hw��B���k	%CD�������e���h�ӏĂ).�ց�%������c�A"j�d;������������/���Ҭie+s%��&y0�M~Gg��(�t"���	�
�r�]������Q8���u��H�Օ�g�3 P����*`C�CO0�1���!J�� {+
Ƶ�/ק�c>��=��Q`]�im�
if���e����vC�
{�#�!e����:P=o3���F˨��[����N`m$�:Y��mB�s69����1F���J���,����i�3����M&��D�.�T oN�4�)�����x �̊a��l��ڴ5��i��\�i{�L���s:[S;�]�+ͫ��;�:�������tW��)�	�̭#S ��"!�%`�q�2�ȸ�
��c�	
H@�W���`�Px1U�����@�HAГ��ab��uwy1&f[f�n7T3�@Gn,C�������=|L���t�1�#�N�G��մ�BR�� p̈�3��.�PTg�Iw՞����x��e�8�_��
W����'(�9̣���x%aױ��۸�[Y&�i�7.֡�YR��#"0JroR���*fR���ˆ�ɒl�"��8�Q�(b��l�t�dQ��E=�1F�� !��CS�#S�8�O������HIsVZ{���S <�uv�bOp�����G&�̓�F1^+����Y�lQqz�§Ma�n����ɠ���(�֖��vpm#�E�7���f��`���P�����	I���f���O?��<^<���Π��m��v���ٮ6qS��瞨�8����% �W�鱬��M�
�>�	��0s����`h5���ړ��n�������0���x�y��o,��}��%��
�λ
N��g�����ð��!c<��$t�L�Pv|mfv��#���;��[����2����=�_��?7V��L�1�H��j �Q�%��l-�3�Ca�'�c-��s�qA���2��}��KQx2�>�J,��|���*+i��/;ڈG�WJP>3o��Cj�gp��#5�T��h{��%��h������*Ih�/��qۓ �@���#r˖��ea)��oX6��+>K�7����I���oAc���:c-�*�����]B��V�4A~���Dڄx]�x^ry�Q�	���h	s|y��c+1�O�x9��l���0K絙Z��%l|Ђ�؞q'3�\ꃳs������̨��MO�<l�Q��i��O�8�k�{��<�Q��Y��nXGn�ԭy`{��V�/diᢴF��Q\0��7Jx�������9U,F�p�׎G[�=J���r]t Cb`��b)�4��D@"^/�2;i���	��"1����̫�j7�f�z�<R� u�2�2 Y�H���$�I�̘�u�Lp�����G�b{Vc�ͼ���D�s�)�zɪ�d]�lV:��;�.s��}h�BFǅ���"o�s�P�@���t��ōK{�& icLѝ�o����9���op�����bbr�¦���FWav��aц#���cZ������^�h��ëD����I1��}<���eN�F�P�?Ce���(�e���4$Z��Vp�h�5r��[��M:���jm��CM�s�s��2�D0Á��=-Y�,�oo��&X=�sv]yi
D��F9Q�5+7�fN��n���rCg{�!����jk�{s���P)W�1����|��Y��C:���G��!�����B�JM��ih��"A�[����
>�H�2�
�kҧ�:�U2Z)�d�a}��
yD��4��uQ]_�Vy/�@#�Z�]{`���ߝ_�D��Y����U��"�`NF7g�ft[ʜ�1|��?�J��s�T��+�e��|�f�b�[�uZ�"��ಈ�Ɂ�a������ӧ�bΝ��+���QQk`6D_��?T�_���SSag|k�H��c+WO��΍E�#A��b,�DDZSڊ�.��P?B.$�����<6�.4�mp�W�.h�����{qa�4R�����h�x�]��"����;t%ΰ�N�9Lݞ�N��8��r+q��5#D�����Wp�x����^QUN��Wo#Ih�	Ӥ0���=�mj�g�qɘ��c��������g�[�o�r�@9�b3`�.
]1n��h�Њ�%���
_�S���v#���1��@-=��o��Et�	~���~�B��}�~�]"�+�EJW7O·�Z�������f�IѨX!�b����

ZG%��l��SګX���N"����r��k,n��/����3��wSZSBm�A�������ю�'�jDkل��cw=*���g7�5�7�E��FbJx�����Nvk#������T���?R�jɔ=��\8�9q���N�R��x�K�F��۵������bO��X��u�w�t�S�Z��Q�G���a�F��|�`����%����SC���螎� ���R�W�q&�m7]��u~�`�UT&rL�l̊�o6�ڎ�,Rdm�9��*?�p�N~K}�Z�ǎ�g�p����}�&)2�ӸE<u0�<���"k������v��)]Tj�F��m�F`�	��DOt(#;o��UP7˕�Z�s��F���Rw�y��>B3��7��&h+0�V��� "�+t^�K�\�����yq3x�x�y��o�v�t��D�3��K�Ǣ(����&�a�.���77?z�ŠT�3x]f�FjQ�q��B6��Zú(�1lǘ��ikC��-��_n�����<W�(��f ��=��N�wWZߤ!M�s6�Ǥ�3�k��3%����qG��'(�09#y�D��^죷�-��5w���<�E-�]@�ta�_����֖��O�W��~�;�Nճ��|��IPL�a��({%��m)���Cb_{�1�\�����d���qy#?Ű%�w^B��,w��-��
i+������~�s���I�Q�-�|�x�e��p.,����K�#{$������W�9��Uw�ts*�PB���������3����}v>�^����1�͸r�ߒ�݅�aY�"�I^F�W�ۋ!K�ٷu彷zP�
�~�J`Lk@�n7!x4:�=�*4_!���[<|qxy�A�5Д�����կ�Ŵ���Ýa �55_ѿ�n�e�^5L�Yv܀@
�.'�=<h�1��^71a�<W��YE��][u	u��\Ϊuz`WIo/([IT:�l�k��9�C��hR�#/]�0���.Ѳ��3�lm����)r��B3�*���򡗂|�+�ޔ�UY��P��I�B���j2��OnAl�W�p>�M�c�f}�	�_���/x����NQ��8{��8Rƪ�ӟ�|y����U �.�~rK��`�_q����Ȋ�7�}�D���o��U~��k��h��d�v���4S
�;.hu��ST�G_�&Pq:8� �C)�0riQ���'���;���t�?vJ4���yQ���ih�`�+��Ҕ/��\-�[QQߛg�:+�Q�:���[���r$=�P�$Y
��?ɤ�A;|���T���jyJ�����!U5�*��Ѥ�k`��s�*��iT7yiD�����o�
��Bb07���0���{��	`ψ�o�{��S��/�}A�3�U13��W�6
h�3�d���<	�8�[3tV��dWf3>���5o�0b>�S+�X��v����<4;u��J+��9EN�bV�'u�Raw���Ȍ�����*�s�h$�G���c)"�;�b+־�KM-sɲH$19��D�}��q*��M)TH
-�6�WZyι�Ў��DzF32~$�y�:��� (�ul~#���x��� 1��u�_	j� {�	vqD`��S`�����j�Փ�������J��R�Ţ���nY��v�iG�Fb���
V�����j�r��=�g�-b�6c_��E��6���J�e�Y����n����tqGg�P�_fɴ��M���ك��:-���M.����?6�b��җ Jg�kh��f�},L|�~�8��%2n�����d�"���}Q�=���qp7�ͮ�#'���ڬx^�F��LI��w(��g5���ff��*�}bF��a���6��F����ۺ+�B��E����O������ٳ�K0Q@ |6�/��Y��(�����h����i7:^5w*p:(��;�es7K����� �ʺ$�~�"N�~�*�9�x膪ŐK=��<|��{)H��ܱ�b^ͺ��-�f^�*��ƈْ��?��e�w��LuI8P�S���H�ld��i-T���WYES6�\9S����Qw�u���@�CIXo�dFlG�En��'@iq��ۏ߮�R	�KT1@.�]�&��Z�*,|n8�����t��;����<�-�N�^���+h�#F���E�tT�3�n�x=��H���{M�/�A�f��P����1G����R+�Q�o�tg�`ȝ�sH�њ�`
9�����9�ߌP?�(����T=��%��8;�ꃒ�Z�i"G�o�\���]�L����,[�F�5�����1�պ�����Ql��s�̈́"���Cq������l�?�K����&n��L0���~XDc)��@ڇ;S$���.2�Ĺ��g�a�F�m�N%�%E���s�"K�T�v��ەq��� 3��hv�2�R��i��{ヹz��~�ms���N_(����z��Y�_ ���[�"h�\���*�a�Cs>���Y��Sk�^��@|�R.�y���0F� g�2Ԡqw~4,T��� �Ls��4#�U�M�,I��v��T�@b(XB��qEf�'Yi�$��ᵟ�\��G����QD}l�ue����
t����`�:��6M�1�n�#�f�q�����N�)����n*�/Լ�� �Ń<��$���C�d�|�rs1a�=D�.�$��ka�l����Y޹x�'K���ktj����R7+{��[sb�lGs�X��xZ��s�H�b�����-E�1[GA<+Ǘ��Bt�(�kJl	p(/�R�����Њ3п.��e� <���Ji��Gw}��Ss����+&E�H�+��{�0���6z܌2�̘����h�w����g�G7�iu� E��&f�>����c( ����
*_Fv��[� �<Ӹ��c����5{��N��,� �����k��AO!��I|�&��t훋2��O
�w�v�{l�!ݓ�m��?.��X����l�K�Hs��r4��+O�l�Ś�fj�Q��K��&mϡ�aR'р 0�H������iͽ�����h{���<��h��:�2��/;^�����"I��8�	��h�u��X�Ә��:"���V��-�C�]�S:���[�@$5�E��B�;�n,��'��9��5�?�eb�b���'�����z]y��m��n��w-Q�՛���-t�Q9n��pJ'�d���r�I�	Rա�^�p��k ��;��tl�A�^����%O@�o��dk�i~Py�����i�5r:ya���]����6�.�&����^�B�!R٢Yl�G���ī��d�g�ѝ�ͷ�a���E�yL#�Z
��LD�@��Hݐ��ة$v�$�]%�8�*9Q5���Hܵ�o �0�akn���E�c��2�L2������8��Y�~�ԭ�>�R�K��\v���:���
fӁ$�^�G?���ɀU���������LLfw�G�J3Q�(<O�#���6`��.*0�ϑ��~�<�'N���
[�����k��زI�=�Ѥ0A�춅EX6�Z�T��{�$ueX���S��*��z���HuDH�Qe��Vc-TU�Rɿ���si���� ��\�;�h9�s@�#�В�hT�T#�!�����~勼n߯]�jS+$�_�A��@Vz���닞Ԩ0�ܥ��x:T��|���$�Ȗ$�3*ic�o}�C��UM � XpT���6��5��*|��wKN��������Zr��\vD3� �_P�&4�v�Мp�kax6V<=f5��l"�0iwq�qL,�0%�1碇|��SiA���g�����^�u���k�V� :�{����L��>�a�G$�K�FR����_�X�¼��,���M7�C4F�.�@��1R疓D�#�Q>�9�#44�����WQ@�_�l2C4� rmx�q��Kv$������/3��<1x��`3xw��0�7� f��M�B=q�؝L5)D9�31bl��z���>����V��y����k���M>v�k,����<()x�3�&U��H,��ݢ9mm�e1.�ʦ�
��}�*!�4�7k<��7�Wl�zA�O��'�X�5�|�n�(���/[�_:!:�!�r�̎��Nv2;���{#'��߅s��i5�X��
�ݭ��p ]1��̺/�a�gv���*Te�i�_/9
�_%:�xۡ�*XL�1�\]�=|5Oү[�_꧛�nW�Teg̳)4St�6�^�Ю�IGQڴjg�{����T���91.r @��l"�>0��lp9�ģ��E�ԉ9�ޅ�5�� �l41�Vt�����bSI��b�PY�v�q �y�'$CƱ�D@Q� 2�A��K}g>��y^_�"�`q�L�9\�4�[�07��R�ȩe�[p����,rM����|Ϗ}��
�e�f�����n����T���2]���;P���>u�t�8�m��kYM��e�Y^vHÇ�u�>+b�G�1��7�� #G�m��K�s>�(Ξ	T��Y!���?oiy��M��kP����9)�8�5entF�1qg"�{�{Y\��=���4Q;f����|�*�(73�S�#�/�=Q�����Y�XQ\��yQ�!���6�<oc;R�R�M8CŜ��oxL�j
��*��W���/�w�cI�Vx�����Ogzƨ2����9tl����%����<��nl��D���V����:+�$b뱏��K��.0I�>��5�袂���>��:�s��zs��U�d�6�g�	7F
Y���x#�h�H��mq�����T�6�_H6�4㤜�ꗛ�)\w��ꅌ�o:������N�괖a %f^Ct��21=�� ��+�Ҵ_mȒ�u�iC�� �+"��e��+�W.�ѐ��pw,Kns���{�,$i3g��:��G���ï�U��"� 8�G�΁���Xm�ɨ$�d�Phlً,vQ͂���L��k��L+�U�Lpצ��5�$owW&������=���&�,xPl�3�A�@�!�gð"��#(J����e7�	us�O������$K���K~̥E�+�G�ןPF.���rg��O��c���;�����|Õ��gN�hғk�%2�# ��n�T�u�Y`5�曟�Qs��~�%5C8M�)����<A�����gP�I]K��χ��d�2	��Qu�p�4�����vPk����R(Mj����z�Jф��a��a�J��k���2��#�Ġ"B��� ��C�����s���>*����.l���2���ؑ������ �Q�/xa�/�v I(��9���Nv�b��._ZQB/�࣎yYrxkK�������ɫ�3V������V��B`�]�FHR��GB���{��^�`�MFK���|�j>T�V��dx�U����M)��=�6�e��]��)^�"��Ye��{&�е¹Iq%���髦0���?�
9��Ņ�I��������R��vh�F-�� �k�0!;�;�DD��F��b�N���¹_�~{�̀}�J��]��E_�P*[n��u�!ԁ�^2��l;��߇���ni6�*�'�����&�,Ղ����x�gI�U%'A��1�A`v���#)�8J%�W��d�.<^���2*{w��c�a��gŖ//?�����%zDW&�R|���,
��^|�l�h�GLJ�W(�(T3���a#��18Ȩh<@��ECž7;�����#_,���
9Sb�y�z%U~��<D+w�V���J�umxAEga9�0ɰRr� ���LJ"�z��3^x&wD��6�zԄ+^m�f���|��aKE���->�g��DL�Dk����>���N������8f�eX��GIθ�\0�J��K�t��������W�}>��BE�M�	ݤ	hΘ��`Z�h�>�;an �zP�
M�Z O�m�(IM�3�~�ԇ�l�9�U}���L���J�+��@5���r`k�g�~PAZV��̃)�V�xxg�Ք
�pR�iء�~���u!�I�2�,R��f�2� x���@���U�ٟ���S��w��Xf���nn��*�Ж���}�#�S����PM����V_u,��|_ߥx�W����K�O���WD�A�'����T$}y�[fQ.�ɩW�=ay>�X�e=�b�.>���u%e��v#CE����`�o_�/p����ۨ"���`�{�B�����O?d�D'�j�}7݈l�)��Yz�Ӧ>����oQ�
��9�#A���fw~F�F`0X�!�W��0%U����ua��aJ�4��Ϣ��[�'����m��������6�;jͯ��#$
)(�R+H���EɁ�d���W~�[!d�U�l/�%~Σ�M�[T|*��.�61��m�S�DO���j?��IA@#���R)OM|�t��{E����bF�{.o�,���1r�?X�G�������5xB2C�mE�`ˁt�{?˚,���+�3;��2�O�+�����Zi�/|�����`�T���A\�Oo�n@Y�$�7ϫ�c�����Xg������õ}7e���H�q��_����R�0Ֆ�%�IB�q֜��D�3�/�\E��<,Z���M~�.�Ќ��m��1Q����~�Jc��9簸.Ӷ�"�l�"��ҥR��Gt G�(v��r����_�8b��dA|SGg���?���HNy5y��q+��k���ۙ����.y{�z�'� ͪ�v��"�ut�*����I�bo�Fd�Ծ�a
���*ߧ=I��H���t�چGrX��^�<����iZ���Nʜ[9{��-���Auۅ׵��;C�T�OV�+����$�:���G��kG�Rx�o/�SN�14߳�3	g�	��r����c��;�o�U�gry���}a�Ok������$~[�ҟ�k,	�Ai�.��`��y\���O��d���=�o9���J����[|�c��䝲�b�\� ��C�Vl�hu��5Ⓐ���;�y����}���f#g �		�ɶ���u�6�&�1�3���=� t�`(u{�lb�g�E���bO����bEq�b2��C2�j���R|� pur���a�h�9�K��9�$-b?M@�I�x�y�U#Yy�oc��~��CA�z�e�Cn)+��G�P���Iw`�M�n!�~����m�R�b��|F�Sa���'J؞c�s�P���R���ۨ���<U%�8�=����WM����]k��O5&j���`��n���xy������ Y�����o��)��ԩ9���m})��r�(�rHj���;]��-Y��;֖o-u�Ɛ���4��j�{��xf;��nO:�{]�Īܧ#��BE2X���NS�=K�K�������K�?lLP
��ӿ���p��22g�;;��fQ�����kZ����e_Q�Q���<�����5�7�A4kv���;
*ʆ ������rY�ǯ��vD-�h(�' �ok��b�Sۃ�|&�(sU��K#SQ���s��@}��'�0��?���ۉY��TT7��?Ŗ�U�݊<n��"'��4c��,G�*f8��CTW�\�j`<C$�kʷ:��2�A@~�t-ŝ>��\��Ц,I6���	�{s.Ԯr�5n	+ى���u�l,����`vgL���+
���&J�}��(S+�"}Wk�(�WV嚱�B��[�c.>�oܐ>���8}U/����͋����Y"[���cK�E%��/ZL�EPw=��Uw���;M��[񤅸O>BN��Oo댉�6~p���J�Я�L=��%�N5|�V��>@ �f3�!�	�xrvv${�֓��u¿�i,a��=��h�2.��0�q֗Ƀm�UpO�5")��b��ٯl��9o��c�/�4$�}�H9��=_L�γ�u!���]3�"Xx�ʯ�O��v<,�
��Հ�}@L-z�3��x���D�aS$�j�H'�v�B�(M��0�()��Bv�Q���+����f=ϸٺ�"��Λ@C�%��{��Ð�ۦe(jA�W��zS^cL8���	�>w���� �v�]���X��p�\e��zkІOd��1޳Ku�W v��ҕ:>s�,4J92LQ]�B���A�;,��k��+�o�!�d�I�$F͕���Z�'��d6U�̝r�R��w��Hr�
W����ill��D5��;w,�� e��^� �Ac��n���T%u$r�9��YY�Bv�+���&����݃'A5�]���ڼ��	_Z����Ə_5�>�����ʬ���ʎ\��
bY����VzV��<=t�%G%�wK6�y!��5h����M�O:i��!�L�����I��P��X=���5x3��ϭבz�������"�5$ڐ_P	I"��0zv~�_\0�?��Q���Ɓ��܈L�=x��x��F���/�V[B�t���ʜ�d~���l0����b�e)g*�r��r�
\Kw�w��]����eE=2�Rף$g�([�ix�@	�;h�B���[>:��ܶ�����D�me��ݲh�}��/�� E���LV�
��,U�� Y^��yo�.����v�EӖ�ճ1ڮV�r�J�:�X}���F~!z�rZ����2KtI�ԣ��^�i�ͫ�(A�/�+�X�=j�P�]��Q.��/ݹ)�hCAc�ÿ�'O���7ꀀ��v���{Q��R����6��&��+9�j�h�Ԡ�0���&�r�_T�9��S.c��Qͩ ���l��_�_�A7Ts�#�G�� k���X;Wk���%X������E�%�+��u���:~��O��ugO�L҂�9F+��E�9�-�E����1pB*���Gr;1{NT���9!���ۥm��>����(�	n��ui��b>��%���|���cW� 1t� Z"qa��A)���τ�t^����R�k\XR��ϝ� �@,��"��u������L�:���;�z�m�vG�A�L�M%��c7RFL������H���~no����Ɖ��Ec17j7=E���ݎ���b��ه�7������gL�c�7��������U"�`��?H�ǕJ�=���0L�ȁE3���_$�K�2l`�N1>y*��)��6>tlw�}�+��2��vAf�r9�j;ΐ��%a"�������SV�h�'�����J"aǻ+���Ղ�ִ��o�6��n�/�"=e�}�)ˑL�5�AC�&{�(�́��-��!���=F��U�J@K�,�A8|�q�hP��\M�)J�W��Y�T�{� s��0�/}p���U��G4m?0�,�i��jmF��J�<�M�	C���v��;r�67���k��ݳJ�]�p�˹T�>\��Y{�A�����j�&\4p������-�#l����w�:�W�V��,�#���~:�12��������n`n�3��V�7D0�,�������"��b�B�0%��|�1��a�d��_�A�k�N���K��`�7�菥iW���T�%�o�)M�3 s;`�T
�r��3�,�*�c�IH�_F{���*�S���F"�E%{�Y�����l����{�Q�5�{��-�S�l]�ɞ�U�S��n�:��+9��2����Y2%?r��H�L\� �]Zv8�y�o�x<0�E�.���ft3�c�f9g��!���^���ʩ���iD�MJTᲝ�K��%̏7�UΈ��'&����D���d�ȁh?^K����VE��7-IK��~r;]��S�
 ��g�hz.����E0,+_���sC�]�����W�j�6�6R�!�L� x���w!�YJ#�2�a(n�(ppV_�&�yE�L(vF�T�[�m��3�!�.Dc	����pE�U����Dz�˱=��t[ޢ��[%���F���8r�3i�r�*�6s�!'�:g3#���&
�D�:PW{a��0m�$���x5���nO��An�r��t�x4u���K)��y{V��n-I�r�Ê�ΰ�҅r�.w����ۋ`R#>���H�����
��2�=-Q��k�Fٌu�S������E݂̺Y+��Ԅ�5�� �U]��w�}!�hDk�O���gaj��ۻ��s�e�=#^m�X!V��ECca����p�]X�{���,�.I��zu�9֚��kN�r!�hl�]'o�|�Ӎ�m�s�o�cvRU�T%������VW�B�w�Z��F�I�6�*���W��;VjE�2�f���|�SOaҥ�ߖ�s�8����G/i�}Y�{�q{Qn�9��؆���T��b��í#�@xݭ�%�F��
���G��]=��w% cZ~��.O� �!�u�����6�6V)1�h��!!J<�x����_z}6#�(�v�al�����s��ܑ�Kݢ���X�sTM�5�h1��t[F�
��\G��L*����֤�ΪԹ�P��
�g�8��Ӥ�*n������J���s�B���A�;^�:$4�ğ�%n�6��6�k�U��w0�����:#!�L'x��j��4���s�>����^!���nI�_ӱ]Ï;P�'!C�#�|�Z1�o����"�Dmb���?;�H��4
����L�ZR{�_iB'`t��5QI���4��k|�>�k���݈%.H	O[(��B���ދGV�s�6г��.����Z�f�k�V���U��M��Ǝq/�K-<�w�X
�A�{;UV�58�ۤr��Y�����b�;<�[���ɜq����M4>ðH�D�VCO{��+Z�Ґ���r��W4�H�Rc���P�:NuXC^��I�Y2�N��
��K.�K̉|���-
H�Aԯ�5\�F�׸QN#� �"��s�;�#������e�dtWc'L��U�jT~�����+�s�f���������a�D�;�2԰9:���W��}��["Yi��,,էmeEk�^M�̓� �� ���y~h�(��^�G�6��2ҟ�r����h���N#�;��#B����hk�N-1���RDF�C��(�*_���>�!n�W6%��-�SϢӥ��f�)\���[�y�<[�^�w-�EY��Z��%���Qf%#���@���*Ћ�_m`� Y=$X���/�t���[�5��w�H�g�ͅ�R�s,�Ai�cqϱ�w5�т\8r�۲���@�W���������X�V��0�:+�@/�G��L}y�����=�܃�ȇ��1��~�Q5^ݗ����}׃�)7,j��2��2�/5����dS�`*S���ɿ�x�2������Yǃl,J�����0������O���ZpdG=��SY�D�=��$�G�޼�y��_0g�F,^nM�Wp������/�C%�59��F�G���p<{ZJ�����[���:z��l��q3P���0s���{�S�ôW'_���o�ZțD&�\)�&�����B�D�@~�-P^�kM�I��ZW��-3�n��Ejv�QTH�N��*���X`��L�MO���y>:w��g�����@!p�L@��������<�m���,���S�g�CӉ��� �.�E���(#������.n�7_ #˻7��Z!��2��`{����^@F����`/�x����gi����W"���͑>{�O���>�?�4X��H~J�_ʪ���76�ʯ���.CM��)̡�'hXp����n,Ƞo�a�;�����`/���Ena���XQ?!�,�Hm'��j��H4y�h�6H�]��Zd�?4�����sp;G<h�E��c��j�M�>�R�渋	q�ݛ�"���F�
���a��0²f��/Ų�{˖���$��@�t���P��'������1<��oT��̈́��,Y�w#�Ӄ��F�H�{-O0��Lu6�W��������,ǩ��k�#�Dt��v8�J���F8��I2s����������0!޶>���_/&w�U"W})s��@�(`R�Uo[��*�+�Oc��p�{�%e�A���� ���y�5��.����r���� ��߫�eh�[���N�Q促)��1��J9�p��z��s��7ֹ��Lޔ�3�YE�߁1D6�.�s�n��I�!u��kk�G��2�e�*�C���U��:+O'�k�%G>�qb�gFzq��lW�N�>8���`8bVXQ��$�ӌ�+SQ�	�<�w$���uy��R�I'(Y���tt��<�C��9�K�`0��i4I��?^����6Q��DQ'��&�i��j8GW�/�眳��ִ��&C�[C�O�JH$=%ۿ*��~>!�l|3�Dѻ�8�R�n�>�_~�����(3�A���o�#��aS�$B���a"D��H=��
���4�7'ߚ�L�J�.�RII�.�X/%��%��B�� ���B���-V+��L�����zǃ��>=O�
c?�RC����_���":
uֶ��Do�Ǣ��D�Ӻ�-d���"��=1��'0�X��^L��m<й�QZr��3G�#S�ݮu��;�K��4�kw|����c��
��0�Ll�EUc�4]9E
YV�G!���h��O��"���;�x�I��2���1çy��2�K�<4ϩ��J6�A_��xF�>�)��3�A��"-4dϰC��T��am8��ׄ�X�$at�>RE�ȥ*q�@eb����C�B<��p��+ ��m|��wcK�V.�w����m�D{��ݙ�A��t?���P3 �Z�Bؙ9�GӍ"���2�	$����c�ܳ�����g����Ӏ`�W��.�7	q�7�#���D���MO�H���\�4��@V���	��؎�g�Ã7�>+�E�e��<�z�\0!/�xZ��EBo�X�U/+rT�#�3exF���h!d�ʑ�H�-��9�jQ��*i��s��y�k���K��Z����U~�8xc��[��Έ
��Fv\�E��5�/:*�Қ/sB�X��A���]	(�~Jej/A ��Z9�O�L!�PC��3Q:e��8E��Ɇ5ϋiF�wD��}����������Y�j�L��<�EUy6�������΢�0{�Ʒ_ˆ"��(�Z�!A]g�YK�?毝{Dy�&!��X����:j:&z����sNټ��k'�b'�%n�
�N��qms���V���1�D5�#u�ːH@9�7��c�Gn]���bBu�q'o��U���K�7���`��7���#ݟQPWMz��oB�H��p����SB>`(l�ET��U��A�����P�6W|G���2�it����v�^x��ǩ?~����쉰��;�e2�p��.�LW����+7-}�~W�Ԅcl[��	m���n>_�d�����߇ޯm���b�4�3'���݊��WVF�Mʹ���������{/�'�2 �5g�cƵ~P�.�h��e��7x�m�'H1�x���wt�R��>���e��<���g��p�Yl���7x��Og�-�C~ ��clB�;׎����8�Ļ�5:�g��E���\�%|HVj�;��f=�	p�.��;E;oV��閈:�������b �'� x^nYP�n^���If�Z�4��![�@�і��Kݱ���i��2�Ao!dr�2��~���.�X�;l� ��6hà���v/ u��>+:��;�F?�P<�����(� ݜ{>�q�ziX;W7�ty�#�=��1i�zU
w����Y���B�&�Xf���)�Q.;@����-���ѪI�2sqd��ؓ��\��n���A���f=&��|a1��ϲ2�8��f܏"�}�@�A�U�	��E��m�޾h⳴=Ł��`�� (��X�N��L�ۀ�d`�l���|������Z����G
�9����i����`�YF$+}b1i�k�S�E�V��b��sX)֚��]�o^�R���L�D���/�ν�.'"a�s~����]�����;/��-P=�΂ris�j�_|`P�%�˗Bmod4��O�s��v�;x�}O���4���I9��+���s^�~�O�,��9@}�s�nKC��d䁟nQ'�8�
g����Z��Vv�x�B�u���<�n���u��@�[��k�Ĝ|��Њ��"���Π����Gũi��K�'&��9��x_�JCFE�̀�< ~�4���J2����|�\�1L�W\���!W���@9���3���ֹz�	Ȫa��C����b�f���Ͳ$�Q;��J�6y�UW�PŇ����~�p5;lQ�����N��X��B V�с����UF�$��e��j��La�8 �5A!g���/�|���T���*np��l̽��`_
gi�~W>M� 04,��^�?L|>����z��c9K�S��Q���=ZK#����%=_	��ѭv�csO6�����aQ��0�*�;E�Z�W�K]6���ތVޗ�u��\�?f]�Q��Ye�)�6k�s�*u�
i��Σ<������48''�? ]�
����'�֪��N��A�3�*���=����%L%<��^1hqiԥ6��Uɖse���N�;�k�����`���!�m\As�+��6��;%&c��r�������W^VƐ�f#5��>���������vD���V�	n��l�
��F����-�������BU-���C��t*&&��a�o���?4� ®����������d}�B�~^<�1H���=������Ų�d2<�~`P������	K.����1�.�3�u����C�б)�	;�\��\���}�h��e�h�5��F��s��7+�7L^U3��,g�l����+w���o��nFS�� �!��9���	Q�ĸ~d��P�e�=�>}C*�d��Ai����� �J�^�9H+�#-T�9&BQ�m��,"o����!ݸ� �2�O�]fSmr+��٭x<Z:�3T�S�x�2�!m�7��M>e~ݦ���:0��4�$4�=X�e��A��������Ǯ����+�|Z��!�z����]}���u�:`T�%ӽg&O��E��&.(�=���!��]8FK�o៶��ψ��ڼ�H���0�t�pS�r�P_�M^��=�;��[�FX5�7�%�c�X�k�~�c[��6F�pS�絍,C�ʝ��o�%�VyGVg�:Q���Ht�cFl?nm�����_�!��Ǎ�1�ga��ui�0�5�k9�Ųߠ��,�Y��q�B��s�2��.8h��N=��{�Z�SB7��7GOx�%�}O���1��y>5YL4B�<��SM�-8t�'Z&m���Fx�6_�c�X�CDO�%����bg��XC���?ٮ��0y������d(�s��Վ�[�'���/ ��0�s�9j��ۋtv ���y����d,�6"���������W��dD$���ʩ��������U�B����m3#rB'��t���bɗ( ���n�$�\f��r|籠� �r��~̑=̉6��?x���nHa�v= 4�*�*Pl���$$�ȍF��<��f⎾Q����m��6�Sڲ��-ʼvAX����T�<3ℓ�T
�=���s��"���I�Ȏ�$}w}��y�;3�缓]�K݈w��]:^��(�D؃O��UBG�'�R~��+�v�x��4��9p��5h�I��l����`���f�5��"g������oF<��P�Ĳ��#�u�ד*镯4oJ��D#L�JB��4d���:[��?�^��*�_Ӧ��6M���4��&����&QzEq�J�G_���u��h@h�|@�ҋ��!3�b�nS�>YT����C�G�1��ۓ5q��'*4��{�q3>H�f���Р/b����)I��e�j��b��=`��-j�]#D23!����e2k*D�+�ܐ��U�y���Y��Y�,9��]����o.J�M."�[���%��|�
H'�AZ�9=�׶��^9tٖ��*ђڹ��	��ǌ��!����t�\�'�����T�wݎ<�-�����1`�mA��8����-a�kA�H>|dWG&�7���2ߴ0>��b�F�+@���|cka��*-$,���<+1* �����j�3	�v�^��,����W�:��ك9)�0"�k�.��W�E:G�&��	�.i�W tvT�J�s�~6o�&���x�r�_��v���f��+��N`�|>J���u�]�֐ ^O�_��f�'�4�]y�ò����q�}ZE�s����H�r��=XL�"�����D�2�H���q��L"�F�v�n.�����e��H.�TX-Zp}u =U!nRJ9]t�'&�e��(�&�d�ݭ�e�^�����˅������F��im!HS�%BP�Z%�Ղ����lF���"�Lf3�[���?	�Wc�dh/Q�Q�A��*�DG4��<��@�㼫���=����W�/�ҽ�,G��Ǌ��NN�Y�e{�"�S����-윷T=[
F��=Z{̴��(�N�$������pP��i�kY���X���_7> ��\���H��㽒/�a��r WL�栥�UѷLn��k� n�@�:�/���^�]>�
e#6\�Z���֐�1dt~ ���ۓ�V�eA���BH��+��v�HJ`!�a����š�%؇�^j|���BZ��u�Qn����.<�m�mIaj2]M)z�c�;L�.���G�r�['���\�Yi�xq�{|#����S���i�����s7r,gw��|��k�(�Mꡚ���Ζ&�0��cInnƤT�?�Gj ؠ�	��b�8�u�C6~�'I�m�5!���4
k�� 9\��~� ���k�l�Q���&@&�%��$N�M����	�1T�rK7��e��S�Ѭd2�&	K9�V{�*H�1�?32k��g���T�c�X���ݗ����G�R�.K��Z�g�&�g��Y8,�)�Ӂ��%��K�a��l>��qQ�Dl���� HA�ra��L���`�4���ֽh����K��1�	YwS��2|�,��^>>�h���h]?9�;�,ֱ�����a�e!�h��l�^��J�UWC 5���_�r���l�"�l���<~` ��c+C�C���Xٟ�R�>��Ka�Z.+������L�����Ǩچ�\�2��U�I*�Fb����w������3>����Po����8�M�Q��N��#oF�v$��sJ��8�F�x�4��4��
vh�����%5�Lr��+
W�Y���6�r}*�u,s��q?�&��d�ٗ���=&k���EԮ�U�>+�b�E�4O�׽W��C@#nI�+�)�@D"�"\�Uf�,���j���6p"���1��H�x�c>q:L ���U�8�J�JV�hn+Ǐ���t���������I�۞ɯ�i����
��g�ʍ�Y�+wݬ*J�+��L9]W���*N��mB֦so�[�q "Q��
I��uݢiC{r��|2. ���<=zxΤ�l��T�1�c����r���=�|�*o	� g6��w2ˎ�Z�_��� Y $!�(��CKSs���4f#W�l����� ���o�}�M�"a�.]��Sڌ/��ύ���4.l�	�����JI�gt��4F>$�N��� c���2���@�(j����H�Z޷�e���~>�s����'{d��R�^���\lŲt��G+�a�(�ݾG,fR胀g��ç5
�,�W�5�=�/�}�1r�Y������C�陫�}� lQQx��08Oܿ���'Ϻ(�1��\T1�*:QJL��*Ԁ��CE&���4�_�O	Iɥ��s��A�V+�\���F�wԵj8eϯ�uX'��B��L(���q@��:��ӆ����a��h�ePP�����/�m�	�"_�읕�!�aE��L��J�u�
���Z\��Rd����ߠL8t�ҠC�=u�q��%��(��!��'���o�.܉Jr�t)*��?�[j�P稹M���{B��]t<|��$���S>��Dqo*`��?�^3�+���`5�X�E[ :	��k�L���g�ꝆS���|����fB�tx�衜�q�!�Z �����e���t����ٸ}};%�k�f��M�d�weu��P���c���s��	�.&��"=����)UJS��	(��kP�HԜ?6�zZ�J.����&����v��X�����	d��#�c*B1q�(X����4Ϡ�wt�3
2�?����}'$t�FVy0ޖ8��>UOU�N˴�<z����%/'+M��;���;��RC� �r|����'��~�=��Z<�ŋu?���xLI�[�Fp^�tP�_�P�7�@`���$��<(ޡ$p�1E9�ژ�GF"hkg��n��y��w�o�#ghWD���90��p�o�����辆�U^��� ���fKW�b5K���+�3�sɗ�G��z�φ���G&R���]S5H�Ɵ��?���F�K��;�˨�Ȑ-"��W��$[EkA:w�4���}����y��g�
��ƒ-�i���)x����b�o����3wT�9����֞{�ˉ���wH
CAٗI|���(�]�� �s򼒉OW��w�)�.<��F��'�vE]��HE/3�)��q�k$�=}7a�S��m�lp���(�W���C�D����W��n��-cGq��^LӜ�qT�`|��#��$��Ӟ�+B6��s$]h����E�!}���<;�����0F�T�I�EA����u�8������@☊�!,_��T����J��x��=1ˏv54�C��`~ph��ǧ�����/K�C��"���K���<�P���j�k�#���~��I��H�fJD�:j��(�b 	YM $om��c5�%��T���%�6�L��H٩O�{�� 
]���U:E�����	/�M�c��$k6EC��a�_e駧z���'a�!��usO���ٻ�:RT� ��yEB�-�Dx[��t�Gx�񞇽�#h��V�8�W���aO�X_�P^ Q�:kf�ah�:��s'��A�:��B���ۋX~=" T��3� o��V~�%J����0M��y�y�-�-�r�mx{t|�]��������q�3��H�:�D��� xr��MΓ�|����TO�;�Rf�p#��U����f��b���T���-�ӔП�����5H�S`��B��F^ƲT?�ѳb���g���:�.J��g����Ѣ�V��FX�X(�s��V����n%Mo���$ԓ�)����Z�ӷ�=�k��sn�������f�7���0F�!D��<Kޙ����*�(�(8�.�V��IoAuL�)&Յ퀄ǃZw�&]o�3�߳�0qh�Օ���X-�"+�M�Cۉ�#���6���{�F���곽jCA2/=cW�dg�������0=|Y_�h��ˉ�f� ~O��̠`Ԏ�3�\��s-%ԏQfd�F��E������=9L� ��Ǳ&���v��-0֦B��?��7��}��/�_��V^�ԪwGRJN�'��Tv�#�B@!�c�Ǽu{D[󊜬�*$�tJ�|����7ڶ�uT	�T�qV�	���o���]B�����n�x�;���"����%9S{jX����
P��;&"(s%%����Q�]��(�,�1.T�ө�?J��g\/�c�챀|��$�k�kP�o��ݢ�a�o��x�Mg7�_�r_�#ȿZ����ߣ�#b�����q�7ٌy����_���r:p1~��MpyS�^=羡�]G��~����?��#�����g[�ƙ�MR] ��M�6�AR�����9o\o��� Y�9��[�5=%�	,]�A��q��}��~k��yͣo�r	�)�M�;�NgX� y�P5�NW�o��
�&��м�ZKd�_�d^M�	Պ ]0�6ǲ��c�=��N��8��)�+���@���UO����܅��;M܆1�{#2��������3��
Fli�S�`Kf�V�S�W�_��[��v�=-k%7�,/�Sܬ���a�B��h��d�E jU`�b��bߟ��(�Q�BQ渤�"�o�4� �U���XO���=7�������k�
#6Y������C5�jɞ)v�J4U�![ڨ嵧(׳�0<�_�������I���>��%cw4Wɺ�䅶��iI�_$��+!�?\�p��ٖ['|��*�bֲ_j��5��*����R#�Q!�g�jT]�4=��02(����J9?�����stvF���	3�Xϳ�)�j���3O�R.�y����rs��N���]��o�$?*͌<&S<��WzI�گi���8$��<�y�r~�»��^ �o_��$���?c�\�?���Jg�V*��.�/��cH�!��}�%�pǧo�Df���RB�8�(}�:���L�,��K58|��bՏ�9o��P�������YBp��i��
*����40_�!S��z�y�53 �{YEHn�˿Wm���
NlV�	���O#��$5Xq�k��2��xI9x� �~�"<X�MPgR T�e�@�Q��O5y���.U��g.��ar�u��&$P�7������z���L&El@�~���?�G������
U���aE]f(
��o8���_�W�eb�W�J6+2T�<@lq�6�K�+�y\Y����5�u�*S��{�o�D�W".�<,㶅���x��e���y�rYl5		�h��-��<BT����ђޞ��Q�=v� 9���Aڠ`� -{������a�	�Q��2~y�E�]	��: n�.P�����h^���O��Z�a&��*��q���+y^'�.��_�d���'��p���S$l�2/[w�c)v}5���Ks�8�$��Mw�0��a�0.,/|����2�T��(]�tU��	��a&��)���� ��E�2�������$�8��sU�T�k��\�z۫��n�Z�����G�m7׿�oMh_��W"��	ً`��� `��̒~�E�?^�Ծ���{�X�H|2�ݚV��'�{b?��sM'\M���E�3t���bd؏/?�|9��|�p;'���;	��."gƑ0dH����`GMlj0]���+��Vc"��KC6��Ȓ�#����FkR	uaAA�m�J��6��}D A�-�����X�����W��S��J6C^�_/��d�����2����ˈ,�#o��t�N���ь�gP�e���f�K���Z�M;_��b����t �h��A��D��O��y�5�J4f�R�J�$҈&�SƉּ)���?��ZM�Xi�-8���b{�d�E���CD��E���YQ#�����)�ҽ�;K���jDX\�;s��
���_�|���?e=��JZ�x�\s3�gX�p�}�,��L,��_��x���R�E�S��txˀ0[�L�<�v�'�쇫s!j�"tǠ���d����>�Qk�'�˻�b�y�#���q�o�G2�]ۓl����#V�D!+�aK�p�XV{�tW0��Wk����_�G��8GYM���PO�KSоH�=��<�S�\��P��C,��S4L-G!Q��i0�<� �e</nM�?y4 �|!S4��_]��Pz�3�rL�w�m�u��.�� �n��w��1�P��/&�i�w��^x�A);���F^2+m����sP5�\��xN�.-�ؠ��$T�h���/ٶ�}EM���bH��cY��ۆ�i�H��(锑�%|��P[�ĕr"�Q>��/9UJ��ݥ�&��,�$!��f�)��"0��.�)D��=4y�B��07�e9��$�V�$��v@�h�ּ�V�,'4J�!�
gD�d�V�x�(��b�Qs��G~D�_�����a���}G��h�dfmaS�V蠃.�A˹,EL��Kh9�����D�j�ڱC�ꭖ(��#��b�E�g�����V��diD�"����i6��?�r���R6�k<c�^Zn�I����	�V8,P��YA]��_�k
�?�q���/2{v�R,>��`H�pvuҳ��*ʯ�Y_R7?ewq���~3w��j�eK�j3�0RBz�
�C��Ln.Fat����v ��,5�ڎc���@2���&Hh���P�6�Zpk,��(�%��n�_��3�u5	(�����\w|��Fn
xEx�Tu�*"�Ź|�y_8FAd�:�#�,+��I>V�B�h Pv�w�G(qP���%$����iL�'�Pp$�@ͷ�� 6evM�mJ��>§��c���3�1�MO^}���1ޠ��:���7��;ظV���I�,..}���w���	4�S��H)	L{�`�7X4����b`t������4�R9�̿�st��:�Hy��c"o8�q&�|��ugG�"Ko^�R���|+%ߧ�B��������0��c9��(:9��q���f��YZ+�D �|�ʣ���{0�n���}�,���Uaɡ�l�N%Ξa��W�p�RŪ�>�
��*��o=9�ƺ�K��M��y�I��y�
p'�F�=3����=��_yFC�F.��1�c��
^���c(�%��_D��^�M�d�%Q�~��9�q�HbY*q�޺�U	�f��+s��`K=*�g"����;��A����P��%`�X#�Aq3���f,�a��@�@xXʌV�1���%#�:у�БK�����$�3cc0�q30�l�3�Fw"�+;ŗ�҆
Y�%����Qy)�qTuS���p��.�Չ�4>��?Uo}�ZJ~�/O��z,��Z�b��'W�Ed "�,΃h��Tȉ�=���)�e���+�1��o�E�`Ihڊ�Bq(�Df,��hQ��y[{�ۤ�q�
���"���TMsh_q�̂�
V�-�"�7�ljY�y�7_��इ*��k��"���s�R4Upt6Ҹo����?���w������i��[I��%�he�(6�u"S�AMlr��ǋs�؍�Z����Ӂ��6��i����X`U<,4��!��`���	���=CENX�Y�H�v8"���v�r�"���!�u����ϯ偪��}��V!�[��N�ў#2�U}�!d���5Rn�G���ڝ$�!��+0؛UIeh}p]c���|��3��:��a,�M�-�wdPۮ-u?:h��؜��'�H�\�Z�#%sU�W8��U�;�u#nl��P��y��4!���J�yt=QJo@�����|�k~�n����?+�d0�������^Dk�/e����΀��&N2_�[���>v��Ԛ'!�PPx]z���a�sk�|T�j|���B���!�K3G��=F���V�)EJ	º�}�A��Ӊ����&j������U�����d�L�:UǓ����&�~����]'6�BS�o�����ب_�˯����ʪ�z��Y��q�MP�~��M�~)*Ԩx�b��Y�'S��չ)b�(Nf0|^"��,h��v+Z��O��g�����b�.����|Ę�n�biHA��hi"~-�y���ߧ���((*�V���^P�dW��5���\�jھUi�$\��m���Y-�$�D�\�o�+���"eG�H��z�TU�������-����B����s��5�H�>s���Ɗ�7趧�[e�LqXH 4%��]�Ty��Z{��� 46=.Uy�o.o����-�r��3�'���au��f�,��>�'ɖn�-̓gx�m��!��>�9�
�n���������}�وR{;�O���'o	���ޱ� �f�T�}�U����<��wDO;�!u��#�Rk�����Q%=���B&/��?�6���A:4y��tUVw	�¾VX5cx��ҍs��I锟-�<���ӌN}׌i��U�\Jiy1�S�3��8)�h�	Rv���������r��FWM��!�A�����\�_t�]��8{BVv�hd�
�88����dk����+�����l��!�YNu�I"UN���Ӽɿ�n��~��s����f�Ղ��w�)>v$B����<h��s5(���f�Gn�E�T_L uX^:r�݄������EŁH+��� ';8�(n���&ϓ�	����2Խm޷�q+5�u�xR�˖�=��B�)��;YŇD�~�3r\�Q�
.f����:�ߑD�#��bZ����Ep>���}�"	X����u=�	B�Ԗ�:L�b�����w+�A*`��*J�����o�y:����ʘ��"d����r���������Z�lY�fn):�N����B>p��v�^s�7� ��V	W��l�
�d�F�곱d�7x�y�f�QU�>������6�g]4K�i�������̥��5�ʶ�"�sg�c�7Yhr��^�|�����C��s?�*b��P�ڪl�׀�d�>TUt��7kyeҟ�a����tp�Z��v�s�BUSQZ����Ӱ��pa�mW ��=u�˨ +�Yц��.)|�NI�˷2  ����1�n|�X��I;gMq G7o��` f:�K ��,.�?�xn�9^����c(���5&.r˰-���ZW Q>�{sr�m�Fk<;a��=�����R"���|��Ī���ץ�"�u��<0�z#�IZ��n����h!Pp�M��p�f�x�4-$@l}mI�H�Q�۩�0q\�@ur�C �lS6�?4��2��1�^!����|6��I��-+�1Ѯ��<؋mbE�sY�xX��K�&rN������%�|�����{ �E��b��ř�NK;�����|�GAzPE�Y�����t�}|��6�+�-1�hk����w�<bݾ��ɔCJ�,:�p�2�i��X�e��ĀJ�\)���6�C�"�{ ����ig�@�Ls�7�] ��e��nO�L�z��u>T��jF�a�4��#ʻ�����S=C�Q��Z`�J��0^+�,�/�"H�����cq��^�U�7̦�&�����yo��TںE�>ּ���|wɏgEZLZ撐k:���|�/.Z��-�{8��o�s��Z�wVfOe��#`JlۃIq)�VQv���zY (jD���|�N&f���w綸�NX�??f���%a=�+Y"w�S�������n���,�ҤR8����k�G2��oފ�y�O[��X�!��Hp�D�6�v�M��ri��2���V{�k5�h&�'=���� �>�4AM�>@�y|�#[oJl`2sT%F�v�!�!�V����d��&[���Y� ��̣��[�uQ�2+@#V��P�1���/�ZO��s�4l��5���ʂ%F��Q0��IXZ_<����`�����m�j�������0|�i�[]w����y�ن����Q��&*�{[��5.���o�k�z�WA����ǯ�W����`^n'mT�)�	��u��C"s��q���3'.��q�I ���vkOV��\��K.����M'P�6	�کW������I�gpѦCf��m|��3�/��}
�~2�z2=�iL�/K���1��a�گ�t55R��Q*��3Ѓ�]�KcDj�#��z	R̯�l�����T��Z;>#0b	ތJ� �u�%��Lt�틴���nj��:�rM� )�e�q��i0��k&�v��� ��[����_��/E�4�P)�|���ov+UX�2L����E1$e]�m.�j�j�(�C33	L��ȩ�(�Kw�)n�Z�.IG
.�TPlj��v��ݜ�E��@�|������E�5l>��i�	O��G�I�)���XA�t'�Ö��$��:+����C$�:{�˹����[��P�E�ٲY����]-v�5�cOt�'/5�=)�|�t��K�p$��m_D�j4��l�p�g&Q�vRh:�����H�-�(ޘ0H썉H9"q���׼���:���<��xo'�?'4��� ���zo���r@���8����?:�s�2<x��i��~P�%<��\�����Ʀ���'x�;���Q[�U�]k<��n �Q1��8^��@+@a��B�c��
��e�~J��)��X��E��D�lqKWڰ�R����M�竦���礪]�Y�5�a!�bc�Ʒ�'�mT���L���X��΋P�J��u�����HVH,�������=�S�~��w�������5%*:��-�6��H��l�M���l�[bpO��B�K0����J��i� {4����bY
���@_�G2ꊿ8� ��\rmkXb�?�HO����i��鈖��	qv��^'�.G�X�QCM�60B�;���f��x��y�xs�����mX��N����	3��&h���&�����o�
� ��Y�E�tZH�%H����k{|��5�[`Jig0��m���|״�p=L�Lj�����<�8\k���v��N���q����b��i��Gf�T I��s*(>���]?m�#���=f����	U:C�қ'���V��_��E�k��x<��!���|=���I����񵸛�;Nذ��?ђ��&pP9ő�/Q�y�K�����K�c@?��`�$ό�������+�h!0)L\ߜ �/BU����5}V��P�=Bi��bu>�6C�ȬO��sIcꕑ �{'��Q�(^!�u3��L7�C��c�S=*�G+��bV���~e6J���|vD�K"r�����Q��T�ſ�hi)m��d)$���������t8�����|�� �iy�(d�/M�xf�I�:WD�3&|�?X$�ywώ��ӥ�:a�7ŷp�b����qC��AEB�bn��0s}d"1BP*	h�(
İ,=C���5�6Kd�7K��4fQ������]�d�m��j���3ׅ��j(��xv� w��y*�U�����Z�쾿>m������+*�=�^V�����<���nJ����"-ޝ���p\�O�������6�l�T�+���X�(�d��~���+�^#�/cp�GA�����:�ɑ��}�Fk[M��%�;���C����hL��N����<(���͎�G+�ER߁���Ƶ+�t��^���.+�/��n���#/Y��@�0Y�k��Xi�Y�����1�&G�^ �@�E�n�W�l/�?�.X� ��ѽ�:z����?�sC��1�ء)�YOtWΊh���-�B��C���)��3�-�pG�钨������;^%�0������{Wއj�]j���S�g�`v���M~�B�l?a�H��Z7�|i�>i-\JO.���vu���t�0� �lW�=3a�$飱��ww�[�eÊ��#�}lhk{N7���>lnOк�^�@��r�)3݊��p%$���ʂ��x���v��4MT-�}�ܣ��E����̑%!<P�>_�EIU5�l���r��,Q�+��C(^��u���3�=��;e
�ʍs�
����"X���9��5%#��Yc�����;��,�SȢ:��5�(�_B���08P�Xl���Ȕ hN�$��˿��ަ��{���U�M��r�?��3��[9}�%D���A5��ƾ�g�͞��J@��h��{��/��c>�\�M#�ӈ��,�64���3�L�ǧ��ؤGT�����t��.�hE���J��tl��;/�3*�z
dO�%���6ٓa�k,��X v�cA��f�qz�}c>���!ks�	��ѭM(t�S3J*��q]��|���3J��B�c��ϰP��S1��d��[��3#�uz.�.�Ѐ #ݬj�e���Ss^gO�O�
qyK-4s?,	>��*�C���j�㡿�i�[)��G��ڣ�,����y4����y4��>?��SY�u>�Lί�L��cȌ|�aH9C��@����R%`|��Kݰi�r�u؋�m
��6�� sS�KF��(V�T��H��82߰?F>���❼l��y�c����A���. H�H��?i#ɠDs��C���l�9�39����Y
���|�+6���"(�I�'�L�E�s�z&S��] �jT5p��u�����:�0G��T�^�����T�������$7��lji��K��nH�c�Gq,�F3I�N�4�U���s����OW*P��f����V�m �t�ɵ����y�4���?�Bw]�����Ǿ��c(Ś��Ѻ@ v>Z��:�.����i;��?iA���W�W�r:��Vrc�d'�E�p���A�T�V���{tu�c��6!�4.~��MV�?�gpX�?��~�G��QcC.L�}�h���9��y
ƀ�9��m9ҸRf�q`�����.T��&�h��i�V|�/�4kgT1�(���V'��f�Pd�5"Iyp ��#�/`Fd:B��=)���op��w��X7CH ������1��)A��p�d#���7=���(eu�Gǔg��~�nd�܊0@�� 	���Y�<7
����Ta9I*Ŏ�CU����HWvt"�ϟJͱ��x���^ �y��9�K����L�&��3��8�	�V�z��rF�^�����u��2���������y��(�b3ӵW
��A�(�ö�8���|�WJǻƳQW���5��I�Z2�qq�-�>� ���3{�Br~�^��Dx�V�6(2�.�	�6�M�|�z�aA_b��,�Î<6>)&�����8��F��^�y?��D��r�'-�n	l� `�1K��������aJ���_P�b���=��k��v�d�j�sZ�rw[
��X���1͕PA��]�$��^f�:�4�߭XO1B�3]AG�زi���j)4�����f�H�͙��:Tz��*Q/,^�}4�����Ja�^pk��������`�j*;�ҚX�aOZ6�2[54*v�Y�
ä�V`!��ܞ㧾��I	�#5�#�'��|��y�9��1M #gԼWh)!0�ㅠeW�8�ַz������7b�����F�L����z�˫gtT�]�C���ĥ�����A���$�Sn= {>���<[�6��r+���Y9q]x�~r�����Y�mV5 �zFRl��Wݿ�3�A�*� ţPڰ��y���k��/������օνpl|�"�Z�P��=�����J���ʂ�vN�܂&�θь���j#��`�6!L�Uq���)������Z��J��j���e���� 	y`B?7���oI�x�7��F�������/�g�{�u����|u= �d���o��E�j�&!?CKb��^�ɫ2��<R����J@7�W�pzǂ������i��f��I����יꝿ�:�tKv�b ���|���2�۬LC��b���4i^��"S�<�x�����>�W!�^ɟ����ӕk��X��E�#c�a�p�k�6�4����E�R�&"H�Kړ,�3:XS��nc��]D	q�6<�˒�p�"�E,E�B�
,_�����,�7f<h�e(�Ъ���g���~P�W�74sV��{ێ�,���d_�r�w�.�<'9�Fɬ<�ˍuJȈ����N��/~�o��	K��l�6�k[K[�����ϱ\��r�n��x�u�*ڶ�j�o���o��I�&�| k
\C��;b��(�	�7Mϑ�(Dvw>rQ�gLA��YK�>a����0w%����X��6��fq<pKޱ,���|�rU(g�, �F&��z����@�N�[�v٧L@���w�huCQ�����w�A���B	x���y���������4�~�E����
Ѧ�F�1=����Jh[�	p�L,�;�F-?v�)�4�vP�]o.ǡd�b�qa���o%��́0K��5���O黼�{��`�� �ݚ�7zWG����H�5"�;a$�4}:�/�v����	M�#���+b���j�8p���KF>��Ũ.i�-7��lw����W�l�r��w���&��5��4Q�m�s���_]�]��$ӯ!o��Ů�N�s�/��&��K�����q��Ȭ<A��F�o����������xR}[����VJ|����4掲��t��6�r$�a�MY��H��m�A4�·@~���)�r �LW*�F����a��9Y(�ٰ�Ma�U�y��+�2ҕN��U�;F���m�Ѧ�z�U�um�!�I�4,�Ɨ���s��A3��%�,��ChD/���'F�*�&�*�u��9�;�.��M��}o��ۍ�}��֋�OU������^Yq����Ҧ�ɸ@P7�puu>���ވ{��`$�2s�{nAvr�+��	ͫ�@�[�������B7Ιܥ+9��B"W��u��(в �V2��К�Gs��

P|�p�S����R���5Y�5�l��,)��SI���VL�.`?�W�2��ف@���;
A��D$�M��t �$������~e���3�0�O
��c���<_��@�),��b7�p@�����Ϫ�2��ڙ>�W�&� �#�읒�|�ȚVMܕ�i��2�n~!���3��92_�e3�7妐FNv)$Ën[HT*P����I��k�1Ձ��`�Ŕ��J8�Z?1t�y�O�]�܂]I��vJS�׊-��s8\�m�8'uV ���%�$"�rWO���V��QCa.f��6�É�I
$��|Z��G�����TX�p#7OB�Ke�s,���n����o��{�p��q�hm�Oe�B�c�B*���ד]�(����7��S!]ȅx���β�Ϲ��O�HP�A�O�OYf.B*8:���r���, �>{:����
���k�k2E8���ߚ�.��Zk���k��U��+������M mюQ�Q� .�X\8�Sk2�枍
���	N�����a���)�����x"�c>.���!��x�0{!VR�����j!F�����L`Hޏ͹�Ԏ+`�I_p����ĥ��:�K^K�Y�G�jy��tF�M��$�J}��s� %���+3��0�4Z��zB�������@��t�M�n@3����j�VVJ%&I�L�]��b�Y�m׿���� N�V�sTTD5ͦ�}�7!%l�׼ޤ��o���pS͑�����~�}6X��(��=r��,��Q�#$�p6|��{����@e:�Qb+�z�n�שd#g��l	$g���<�?�� τo$Z����'�/�#��T��k�&W�a�`�5J�)T�Ps�_��&���
�0����u�  �:D�-2!����㸻��k@6jq��|*�����ַ��z�{^��!G���
�'����?d��)� ��4����
�Osu�;���B�*�J��e/�j�ɮd��<S�^슝'4B���, b���	��u ��s)l��j_~A��W�}K&~$��5�C���a�������b�E�4������À�ED���I ���Ŧ�$|�����J�����t�M|��Gx�Q���O��,��B�OyʭL��fiҏ����ʗ�j�Y�0
!?;�tfv��)1H)��溭4{f����B��\�-T1��/�:�S֤9�U�36�Sˊ�7�-�Y$�s���F�*��^E�F�h	���z��yΩ��x�A�%?gvms}x��Z��V���|�ƩNȉ1d��DF��劗�g�A،a�	)iɨ�����0���s(��g��v���,*(�~��k�t����F���
��K��"���t�ɒ��٨����zp�o�����≹<���Ha� �	'���k0�R������+�;k���$+GxSbkF���;%^X����r�T��]�j�,α7�!y��2oA�x-6�Uލ��0���d���Eѻ�<�Ρ�+?3N�s��,�X~1W�O���#7QG�8������\���snE�tY2yT>�ߩ&Q@��P_�T�|��^����fp1+�R�<�K)�q�꒒*v{�a��Z�D����S�DA�����o�$�6ڪ��S��y���6�L�gd?���=6
��'��;�"J��ͅB�kr<�t���Ӊ)6>�$��^5���k�j%;L���p"���F ��X�%*�Qw���fm� KzD�Gp����`	��8�v�Ծ�!�a��Am�!��b�ɚ���h��9 [��9i���h�>�:3s�joT��z��e6pB[C�j<D$Z��[n.��
V�F�60����y��2MN��r�3#i�a.S��Vz��_�'N�N5�\�SNÆ��L�i�V�,��C�/(."`Bit�u��	v��}�R�[��>�Y�A�f�*}�|)�4r{�s�!5�&��i����}�
��q��n��.Hr*LP�Gͮ��� �K�yx�c/�wK�s�ƛ7��EW�+v~X5��*�Φ�E`�V^I�uAGǎ�ǿ`��jA��cpM˖<u"4�'�iK�U&9}��aN�����f0fѻ)����3�_[�:�.q�nM�5踧�~�p�7�((��zП]������%�mQx��t�N��4�0åJ�������E�b�,�x`("�LWX}��Q(��V�����m�9j1������Qc�^o�S޾����.?�5u�W�0��!�4a����ρGߺL �4b�> �0�s�D��֏�ޏ��Nd�>I�3bͮn�׭-WI�o�O���;�Ƒ�E�!Q�V����
��/>���.&�,�Ċ9�L� 6����L��K>��X3~-j[��Ԥ7P�B��I�H����+Y��k��?�J�ԕ�[�ixؑ�#� Ou���m����ۤ�$�$��j���[��=a��B��S��aoP�g��&�̰[Eө8(3s<#W�Q�Ɍg�<�A��?]&���R�eUޢ��xXAU@:M��	04g�W�����'
Vك�/69����f��&�=4����d�x1���*;�tXL��2A�p�8\�.0S�"�~���U����mvHb0��zi�%"�i�(�F�i.��l�s�]WbìL��1}�,��oٛ��	�2��VY�����^�� �?;�7X�����%�G&F}���Bd�Bc��|0���ce��<����}���d�����JQ���tb��A�\�g�G�FV3��V1���U;��'�r`��k<�r<��O������E��;���neL$��noϯD��	����K����O�=-�01(Q�y+��m�f�,�	�i^,0�Y5y+�+0}��47<�������ip2ʱ��|�F*�_�7iT�'�Ԟ�u�;޹���<� ��X}����Kܑ�V�a�L��a��~K���� �:%���TW ��1�~$�߯`�߀ʤ�m�qy��<$�9�r�:�{�\�fZ�/B^yG�*��&n�(|w�$����qԝ�|�mm��i�Q1��)�%�ֽP�Gn�9�PO˷9��C �E���	��Ӵ�Щ(E�A����:�9|�	�o��J������^�QKⰩ9|�4��q����B�M��j�0��I���õ�:dA8�|׭h�$H�E���Ap�v/%�4��}~�3��?GX�Ƌ�";_�U�=Xٍt��%k�φ�>��^-p���g4���;��v���r�d#D;P5w��j��`�K���pC��b�E���їF���:I ������������"�h:���Vɷ�A�n5ЕFh 	=5��sA6�qP�蛃Et�L��Bi��9�x�#VJ^q`���Eb���J�l��Q|yҌ!uІ�Y�2��`������zg><f(J�h��-���cr��^#�C��	�N{*c�V������\-Gھc��.�c64{�j�1�]{p<-o�O��Y��c)�I��� ������Y��13FUF�T�2��C�I�a=u�]H^[�ذı� �l3���hG�+�� ��+���"A���Nz#B嚞p ��z��-�6�X��ϻ`��5���?o>�f� b�;��}d����V��s�v
OV� �}�*���# '�
�z����,�H#녖�J
L���I',�0f��N��n�%${�m���OR�U�2�S�tI�fn�+aùE��k<��D<@JjU|����(�m�ݼ3�]ٴ-����OS7_U0Z����ps��s�t��=���X[n��s\�t�Qs#����p��x�nVO㥑;VK��-G�ck�Bf�b�s��ͨI���J_�5C
(�0��G��w�I�����H���	��!Ƣ�;cu�0+�\�Q��]�'0�2/�jȵt��!��$N�ν�