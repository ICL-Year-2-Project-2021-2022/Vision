��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P3K��$�?~������\͡��dk�⍥xm3T��8�׬����:@Ӻ�n~��6�*ݚ������a4�**�1'wO���?�N38W�'�T�u/���~Wpm�ك>.��0#�����Kj�l�Q�Zj����_`�n}�T~�w� ��v��x�m6�f����|2*��Q��^�Wh���	3�m(uuc����h�K	u���@��҂����+��=}���J���0����}(U�%�c�I���w�$���+� ^z�e�kh����v|b�>p�|���;B�-T|�M�AH�iUuN��%��'dyHpf�NC����r�5@*�T������D�ʂ
$�гd�S��zǕS��)|X?&���Z����N<e�uQ�I��\�X%I�LRj���-|�Ľ��(Z�Ӹ*��9,.��d��&Q��ǀ̾�VR�4��O�t��?*�E�:%m�v�AV��t{��ۦ�Vi`M͌y$��o��K�o��AF���59m�Έ�N;)�c��MNL����U5��?�����c�V�O��o����#�E�e3�hBƻ����(+��Ƚ�/���vQ��G��`t�M���&��O����T��1NOٲ��A�N��! �ozB���_�\��Z�w�蝀�5�G�K��K��߸��9��~�Й�`w!͇��������b��Z����'S,k�l�tȱŕ0�y]p�U���rE��\G�k��=�����!JziAϽ"&�B9c�ǿ�� �<������l�T���uO�L�G��S_n��;֏��ݻ?`w��/�qH�S>�O���V����K3wv�
Z%�:��o5��3|�S�h����N�u����Ms۱�b�m1�;ewiXX���f�ٺ�w4����*A0���*����g�����g|Ϛ�چ~�r�懡�$6���"��),飶g��n�V�#PVg���`��'�O����&H_򐅞��U6��%ܥ���I]�t�d���W�&		���sSr��`8N��`:�"[V8א�3�)M��!	ŷs+���|=q���ɓ~f���4����2l����k5�e*��X�l��Qw c� ~���[�A
-��O2���kW@���aj�~-9�K.���QN�Z����%�}�5��mg���a�T��fV(q�e�e��L݌̯�|]�^�K2�O�v
�_Tg�����)�3J1��G������_���?j�Za�����@�&�A�ưKA���~/�/��0`"F��Wz_���s�ȌDAK/��GE=���q�Y;sǫ׸���s�!,�����`i�z�ˆ��"��wm����	�:�#ho��9��`�Q����b��+�e�O�ܩb)�������m��1��G5�����8tN_��q�[�����`���p�H��}q>�ʠcM����+ظP���$:��kȫU68A���6���'��}����ߖ��J����w<��>F���HI��tae���$�J����*���]��|�E^�3Rby�;�KU�T�s͡�T~��(<Ϊd6��Ύ=AZ���� ^������F������e�u��?��M
��`���cn� �EF�x]����.�`��U©�F^��z2	"%������6���'h���WU������+�9��{螹������;��HGW�4��mR)d��c�i�δ�9��̩����uF���;8�y���U���M�O�+kW��>���_C����O`�� ���{�}�����{�N�xf#�&"C#�Z^��t�{���MI�e��A_��AJ����-q�"��R8�ܪ]_�`R�?H}�j����v���%���6� 5HM�$�#;iw�5S'��uhywȎI���V�XFc[|/��U������x�.f}�]��:�M�dn��B�6�v����E�W�l�2���F��*#\�%��`�x�(��17z����J�p��>�Q���م�����n�a�k.QޘF�qay,�������e)��#����r�Sdy2�h�c�����DD^�@�	�$:�ôX[^;��~<�6��(
�����u�/���{�� ������P�fW��;h�����뢢"J�S�#bh�X F>��n��|2��fN��~�uki2�����H�1��[C�3����'��ܞ|��W�4[n���������{Y���6�5�g���d;����x�+q�(�f::��?\lF�P��Y*A�w��Ȋ	��4RG%����W���%�}X��Χ��70��]/��xr���޴Է�{>�-~��b�ë�9� ��=�x�%)ţ���Y�w�-L����҈'`1�Mf2�(��?�R�?�`BN�KD���'xK�,V�s!�x�1l�J ���Tk|�hc�		�H�m!��Ho+�9����C��������$Q��{�AP:M,`����ekZ�$w�E�tF3+޷�l����uE��fQ7�]e���}+����	C�t����Lj��P�\���U=j��j��3t5%�'?�>b�5@}2d�r�Y6d0��\n5�,���݈%��>GÃ�N���?�R$%��$����B�&�ŎҦ��7?�|��]�&� ���_����s"�ssI���yP��.�>�ŷ�=�����2'6�%<�����̕ #�'�5����* h�I�������!w�ANb�t�U�Oş�0����]�0pf���l¦Ŏ��_�Uy��`oY�+��M�Va������9h:�f�����*��Ѣ�$}�:���{�@�\NjA��48��
��ڥj��])� �)*�݄�� ]�����g#���oL���a��:�j��G,J�{̖��ݐX)΍,���j#Ia5��%�W�r37Q��o�QF̵��%�q���4w�	�^ā����א�S���8�Ť��d6�~��M�9.؉͕�hk�+������ ���8��=�Q� 2��n����rŕ=���{�9���3�(˴�o� |x��|SKܗo0�o{���>��h�p���%���i<nX؟2ͣ�j0�}U����@�g̛�P �/�咦���>E��;	b��eC��֨qXJa�cS���/HX�� �qse��2cu1�2��4�Y'Ú�	��9� �~���ZfY	�7�%G���u��9=���F[��^����.��{�('�J]����S�������X	��l���k�ӽ���|i��f�~c�p�ȒΘ��H�M����
�"���*r�((3�b!
 W��_�����5�!-�Ϧ)H[�tqRO���q�m�4 �U�ȇE�;����L�c!�QF�_�鮃B3������6!VPN�ɯ�k�J��r�m4q�>7�[˓�����]8��I~&��l*�5�i˧�8�.M5ԉ�B���;��^�u�1Mʶ����0�K��*�}����"[k�B�[�s���V;-��󍯓� ��7Q}b�S����	b��?t�^����;���:Yr�	���:Lx.mh,;yf�gJ����s$)&�<fZ�a%+'j�_��M�#	��T뻜�:�т���Y���=��ۀ��P�J�Y!�Q�JJ{,�^��`��/�z,�U5��+=2i��2jn��5(l��Қ5y��r�_���iP�}7��^��o�L̝A��v��|~)��b #���"ϖ��P�e�4�9�A�#��l`�Ėela��
*��9|��ɲ���)���c��8��?53�v�������`i;��Yi^Y&6jg͞��7ak���S��ztr����b���o�Ys�B����4��d8@�(��M�4��y+ԯ��
Q�kiۮ��!ԜbGtگ��ڥ��Ѣ��F
O�VD�~�9���,������Ő}O�C����i�x|�HB��Ý�[�א�f�*�\��EC�ec�Վf�/��8Z�*�ϛ=���1���S8th�]�w��5���>�����2�&�iӵ̋F0���;�h�:��g��_�Fz�^&�!^k�@cQV�H�����u�v�om]�0�˾t��w��R̡��d)Y�7sfn�v��׎���z�H|z��@�a������Ó-12D�m<�!���Ԡ�t���e�Sl��B���l�ǃ�.|��W�Ɨ0�	=�����|�@K�Ae�������y��T��Q��v $��l�2ڙ����vj����JRdX������,eM���}��/�/H���j*��u����Z��|�ņ�ID�ȴ@C��Ӭ::�fG{�X�����8��mC�;L�[Rސ��D�/�9���e<6�3���j(l(��K��P��ƺ���������I��F�0Kh�7�T��&.X��Ei����v,'Y"�q���G!͊{:���������k��	��<����_�!~w�6�o�dnxL���A����S�o�s_�G�i;ɍ��q1d`A�=�-z��J�I	�V���j�I���y���JV�
�Od#�����t�����szd�i��y�?����H�6����-ts��V�6[��Kj�ΪWhQ"��Ak�<��=R�`�&�G��{:�rth�ꮠ'�=M�����mp�=��T}������`�x��RŃ�E�m�$����_�/AK��A��'6)��N�]i9/7͇�E��������aT��ԯ}�F�B��R��9�+��K=�h=X����u7��H$��S-�	YL�OZ�Jvv��_y���oj�{�a0�*{��H��r��?p�'��ġ>�!}�z'�/2U3���h�5��_$:��#ji�#�o�D��C��TN���J��|V�Y�0�3c�y�K��O�J@������D�Su*�{r�����0`[����v��=t���=^:|���
XL�h$i�@S����ZT������S�=BŃ�َ1äKh��И�c�9)C$CI*;�@N�  I$]Go��:���tQ�.�{p\vz��0�J���w�fv��	��!��� �p��K��96*\���<�כ�W6�d�U60� ��(l�v@�\��˩��τ&�H�t��%N:��w	��2�M,�C���b��G�5�I�5���ί�5R6�"�g�c����֑�6��-�Z���
�@(ّ�<�L3�����J}� ߰L�*���W�+��6�&��ي�E��T܂a��T�@>F�>�Q�I�!n����Ј����敱u�Q������r��~��s���	>j[�{.��R1aQ����P�NT�x��,	Z���}�eq������H+�A������j�e=�j�)]s�� a��*�t���mE���um�b�J�;fc���8b���s��s�\Zyk�f ��gWO���W���@��.����}�ALʰ�tE�8Y�DɲǇ8���w��G^�E��> n,���c�>�Ss����EDO��������(�����S{���tʨx���/��+0�P��V��zu�'m���-}m�L����DB����k�%��I��������b"��&��V���7�I7~�z�{oG�%r�"��KS�L�Vt�L�����y���Q;���4X�c0�{����Xt��NQ'�Fk��^[VC��[��X�Q4E��+}0��;Si�M��`4Dj����5<yŎ"J�>6.�Z9z�ɓ#L�=I�q�Ո�H�TC���+Q6�B�r��a�u����|����³/��2�[K(ڨRj�"�$�����L�j�[�!~!'�C(u��~6���'
n�H���\��k�

���HH�]�:�6�(�71�X��yt�&m3i��FR!��/=-k���<�@o�Č�w->�7�݂ױ�	�°���K}w��}U��b���O�˹W�y��`21��hm#I�8�Ծ~�sE�h��T�	���s�?��~#��k�FV�&�܉�I���A7J����=x�l�8F�&����dY?���2a$�[Z��Oef9qI;��Od;�	k�)5��3lw�Z�#�ÐǏ��W��3������|�����=0���J�v�/�k��+��qS�C�`t�ޣ�Ӡ���ۖ<�ˈf���6��I������y�,��l�)i��܌��t8Z���k�qm$��M�yTW�xOO�~#N�P�ٵ� ٝ�巊͜�Q$��:��e,�m(_�%9��ա{����2c�)Ŵ�1q#�c[s�٠Y2n������ҙ˷�2லxQ�[wMa ���i����1��ܽ��a�
:�\�ќ�1h�ض���w#�P{x�^ճpL��c+��+�RΙ���j�0sT��K����@T���<�|�-pz�[��uO\*z�MD7v֞�C�ߡWXG��b��p����x1J�	�19VӬ�"퐨{I5u�I��k�s�8q��L��;N�4�v������>����K�Z.?:�����䯉��~$�F�t'(-v�E�-G�9�m����n݇W����ʁ�Y5���<L"���#b*T��ań�k��_��A���A�ΐ������j��QⶬG��Mp�cY�N'%�k}�mW����i7������N<�L��S�]�cf�u��h�,V�������'��[�L��+P����Ȉ4uE�{8w�d���M�ܽ
Vޤ��q1z`�%�g�h��� �Ժ!*���*E���0�ήp!��af��[��'l�+,"��7;�q�����F���lN���KZ�E`^˟~��ƔG���JƺE �7�0�u�n��nxZ%�}�ෟ��m:b��@��[ ����\��uo��X��i>H|*�ZC������4w�S��s������0�W&ܔZ5-&We�	A����N�:nY��RɉJ�5w��g�Fty�c���/d���b@TL+��oy�m�8��th��Cq�,�$x�̒q�kU�Ȱ�H-�%Q2��X;��	V18y�O&Ӂ�[h��,)�I9�:-;]�+����i�/7걀[����aI�뿇�!�E�
��P�ը�+r�)�ҝj�����"'�������2�
 ���Fe7��ܪ&���0����a���)����V��*�ò��p�u,o��f�1gd�U�|��_���&yǑ��Ymzc�2����j�Y��u���siPH���렷��"Qǳ�[�%m��@eƨ+O�Y.m؊^���0�zP��u�Λ�l�9��(����3^J�WAt]��vfE�`"
f~�hO��}�����K��,U���K���6��s��TFsi�x��R�#��h�!�$��-{�� CG~%�"�THnǝC�� 0{i�ď����`��h,�^�l^2'�YT@��"��7F���
i ��T�;��q�̻��Y%�^���ZcW�:+�܅�<	9���T������uJ7�ـ�� �_���G�o��{28��5P�'ch��F���⏬�/��&ժT>0ݦ�7�����qUx��=t�/BozdO�@s���Q���NK(JθԉML[�G��?C5YT���^S��k��4��aC캀H[�)���e�ͨǹ�z��
sbf�e��m����Ĭ|Y~k�����-�D���߉�3�2�P�`�+���d��ع]�*V��b�������7��h�ݵ�����Q�����-�s���
�lbN�=��Sܩ5fŕ!��@m!����\3���2�V��Q/��@�M-	�� |\��}�9d�Z�]���_�p��v~��❘�n7��Z�>\��%�&2m�Ƿ��]���ƿzE!̆sQl�"�i��v���k��,���TQi�:�M�F
Ű��=g(_T$�"L�x��0Ō�?Vs��
䐝{����k-M�5d\��d�i}*�3d�Xw�w�������o|C�3T?�3�����Ԙ��P�,[��v?t�a�
��$��Y>^�`������]e��/����)`l�!Q����3�*ب. aP�����2�9b�L��fBre?I�W�"�K���s:����(K��t�e�������]�����ba2)|&����4x: [n_N�&R\p�e�,4�U��[�S�h��M0��u(��g�+�Yע�k�����De�V��f���?�q��EZ�Z�yw�Oٸ!@cW�e�u����	�()'���
w�F�7�(x��y�$59�JF��I�jG;���$dJ(|�\�WB0��A_�Gk�K�,6
���в�L��׬�pO�N��ӎ_�A��-଒�̪��4�U�2��X�+J�p桎����dH{�Ʊ=��5!�@�7eY!�}`Rԓ�.s�f>��+�HUKB���_��yܒ���<��4�ӣ��ċ=��>XD��뺸$\j���m�諫� �>�|���.��a56H\��GC�Af6�%����ƓU1�I�k�������桏�__��ʺ�f�e­����?�>���\bY�k���Á�P���R�~[J�j"zXR�b������߅ĭ?	�k�?�-�M�;[�����$��ZX6�����GvqmPUc��l�~j�6�i�̢&����^�7��=�dc�m
n ϲZ���]IK]����RR�;~�˃�K��q ���)*�*n}���O>�����0��E�QM4��0�{�P�(���n�����He��Hόr}��#���:n	��xŤzê��j-A!�UVע�5w�ׇ��0�}�����5���g��<��9b{y���B$�܈����b򂸸�{d�, �*���7 Ձ�gU=�qX� ��?�������G������}~��-�Hd�i�4�qq�U��
s�k�s����
*����p���a������"�Ε�2Iŝ����&�L��lG�]�XU�=��, -���M���Z�9��K�P\��A��Ej�;]����VbP������#u��Oi��B�Yy�X�`�����]-Hf���O^�Ұ�E�i�y���O���;�:�fzI�y�&�n��̇��gu��\�M����Н����j��r��+]XN,�X�@�G(�2����i�~*+��s�AU�h����
�=����	2�]@Z��H���2��ʏJ�G��]�� �vL�=j$��zJ�6��H4Qկ��Ũ���(����-�J�~iW��t�Q�	E���E�倄1!���v�V[�Eܳ��44�2��|�%�k�`ǧ�p"h�pYn�z�.O�*�i_��0��7;��9xЗ���.dz�9���F��N	|�24Ǽ���G��ᵀhW2���یH�E�mP��&}�μ�����w����Ymi
�{��Zۛ�ᮐk�ˤO L�B�{a����K|Ӫ:�N�̤+`��,�oXY�SDh�E�������)r�9ƻ�_�_.��0/M���Do
U���ź�k3����Y<������L�z�,�3FD�&S���V)>����E�	β#��L�ϸ���1~�3�gߞ�,�gk�&)S�p������䏳��3���J6�b�N����$���g0�A�����`ˁ����cVi,%u�.\Bx�T�P�k]��t�����Т�i��MzQ�3[$���Q�?ZR���/j��MB��U즿���[D��Q�V[�S׍���/�,����޴g���(�R�`Ti��Dj����mO��n�Ў�J�mߖ��z_�T�4b@:+�<8�I���#L���
�"ް ��<��Z���
��ӌ��x>��w��_�ӡB�æm�Bi������h�{�t[�3?g-��L�?�Yf*�r1>d��\=[J��_)*��.�����3yQQ�4�O'-��`_��x��(�-/^^\ �c���I,DTG8W�ꇧ�vE/ a�D�2���]^&��Ӊ��yP�5��z �W��^�8ɖ���$��Q#>��B�v�5�q���������{���V��ٸY�����V�@E�u����T�i5fre<�1�:��
�_sC�I��6�~&6�����G�=�%�V2)���P��yqZ���<��W��8�z*o�*O���.���3���ő�]��OMħ��=v���И3᩸�f���w,  �@c�=ҽ���Vy���rȀK!��b���a�TGn���.�_Z�"=l[�H��7�̾��^�C=��c	*|{�<O�j�C��v�F=����:�Z����`/'0���@GZw�d$������&��cJ�h!@���Dr8��}�n��¡M"񃯐/LЍqksএ種�D���\�|�����Fu{V�HCj�!���p�Bz�(L�#ʢbj*�����m��x�X��9��u�����?��>aH]ʚ�}�}���ǘ[�B�1:��`r��_���騏%�����@/ѳ��MR���&�0WҴ� ����}1�/��ַ���|��3ɥ��4��*�*���o�"���ۑ�����s������g�[b����%�f����j̲U�-���/��oc��t����%c�����L�>��s�TI.�/�L%�Mm|�B7�_~�}l$����l�A��� Z�$��m$�
�D���e#^�C(R��|u8i��3(�NN;��A�z%�	�ă'no
�'l~�:o�p���YⲮK�GojN�@VgQ��Y�2���V[P	ա�<�{K�=N�.ً0?�
~m+F��0�F��u���<'��y��t�(�a����7��֤y�9}�j�C�ĺצ�I���z�T��g�����Y���j+��5j[�fss�ǣo�㝾܆ c�@�N�!NKo�7��ԛ���YG1��{˪x��R}r��@�D�:���Ƀ�}_]Њ�X�پ�rx�E��Zﶤ~������nϰ��+�`��<��9ķ���ʞ)��]��x�N{��<�*�6p�<JZ+'21|s�$a�W`h3��R�!!ɾ?�^H���j�|�L��]u� ���pbQ�����T�Z�4�F/?%��F��H���t$h�-9z"a�F ����J�kZr�闢�:�=�/#:�$�0�a{���(}�Ӓ��a��Sj��(�%�t�XB�������G�Qc��aL�D��-�Ƴ��uL�|\3���k�/���%u���H�(w�5Ah[]�Oש.ҭJ�kp!�>�G����2PT!���r؊"�B�pϡ��E�G�3���y����k�(m8����*�<�s�6;�%U* LHXd���Μh{�
kX:(FpU�yR�6��g`d{��8�dpʗ���4�U�iIK�lN`fM	� $�/׳��ql�a� Ub��u���&�
�3Z�vap؃�?��o���t�B:W6l����:���fM�ň��	������5%e9�V`_������N�ȸ������ҁp�~��4�@�ӯ��|X]Cct���s��/�_���*��]-�Պ2O�����"��u_�W�\�
8�u+����sA�?d�;�"�y|W�3җ���@8]�w�[)���b�O�,d|-r.qg9%����l��{�.[c�I�	�0��Dm{���#�F��b����?��tG�z(&9ـ�B z+�UV�.����bRU���E�/��
a��j~� $3�>Ʊ�X��ߛ����1-~�:�^��Ї��'ǩ1N��V���"�{��7)��:Q�`WT���_I�!�2�Xsֱ<�b�70+�$�$�K�����$��z�)'I� ��|�ADRjs�������	4w�Wi8�����~IQ8�>5TmJ<Q��sƍ���%f	��M�<%,ɓݷ��7�]1JX�hu-wp��
l�'֧��-\������6;��.iM|��33��LMj3�:�z�+^I�yg�j~���zz��|LK2��׻��$~�b��M�4�to���؉�n[h�b��ۖd�!�`����H�̒�īG6Lզ����cl�8��U��,7o�آ���k l��4��3�
��䔕P�?��z��+�/u(:��C0[�c�n����H���@�̶�h����a���k�C�q����k�r63�K���71���:U���T��[�P3NeQ��m���%Q�u"��*�j]z3Ʋ��������ܘ�����e�)+M��b��㏧Il+j���{��Ɛ�v�Ӛ�vl(cV����J-\�� ���ל�/������$CO?�>'���1�M��~�#�%Ge8�C��t%;�8�c���}k]�xN�h�zgBQ:��8��4U��^Պʻ��R�����Xȅ4ŷ�F�^���J�_��?Q3a���o�!9�s�h��,�bM��dE��>Zx����xEv�y貮�EIjY����C(���gY�5N$��fp�/��s�)l
�#MѶÇ�bN�\�ӻ���
'���#�~fD��p�Kh��t��������dph�D�D�uq��E�q��x��H���YT-F�����H�d�W[)ci�xj�X�ޛ����7ȂL:p3�]���s5�)ɀ9�S�N|�����
YQz��憫��& !��Ķ�����B����u~�"��u�x.��3}���D���{H n3�sH��"OD�����siYW��P�+�Ij����r��1�U�^��?ް�θ��' `�F��!*q����{<����8V�2Ɖf8<��?������{���O�ko5N�8D�1eQ\fr��Jf�fo-�A_�/^�{��܂j���7�gj�^��R鿟�󙪡�y&��s�D����O���.�2pM�̫�!���yG�81Uy=�h����O� K�bw��� ����L���!�x�k[?բu)�D�P�{h�Ї�����&��8���#�g�ܦ��O���j{�}Y� ��'��ǐ�E �ē:��(h�p��!���l�dM�Fx�b�5K�y��IZ��U�B�f��mp�Rq��}M�<�\
�<�K;�&������L9���PcU�f�5(b̨�㼯]��!�o=B��1 P��ϱ"�哦���'����M)ϯ�<T{}4)�+��+`�\��-�;�a��2�ƈK��	5�*��F%��L�d]���U"a�%���fq�S`5�W^��2e�
����O� #Sk��0�y8�\XL�?7���<������i:�}Q�6�+T	!p�\t@��k>%U�MM��ʟ�[KθRx]�+�^�Xw䄖b�9����z���+�[e�SGG  V�^J~�M�ȍ?X���u�n%>�h�wH+K��C����vڱ��{� �{l��AzVP� C�0C��[(�>����]'�}d7$TIǁ��fJ7~�S6��Kڑ�!�g?P��ltf\���Q�����@�h��Y*�J6��3'�I����^�FL5�J�V�i�!�H��U��Y)��3��>A��3�5�n+)�i�o�r'�������3?�fĊ����f�\�~؄_Y�*@�" ��������Oy~ϔ���*]`�dW��h���/]�:�5C0�/�&��4� t�O�g��!�����y���D0d_�IX	'�W�R�*]gRÐ(��&�2'˒\ȩ������&0$�[Kyn�;)��%Br�"�" 3 \�+����Dg\|���S�M.����vk�\���A��0����5��n��.J��m��vx��ͼy���9��;$5M%�*��������R�"�Z{+龱�����9������F2��*��1~ ��9�:��/��F����<V4m�0�-{���ض�z��sbfa�����Խ(8e�̅���W�1PzM�;>hn^�(R_��ߓ_���rA��g�*��VΫ� ;����w=#�>�=7�uu7-�/���.&*�oL��?����+�ӂ�W�x�_
�y�FBG_|}���Z)���������Z�鶾��>l�-�<퉚3?슧�3s
^��e��U��7��q����dۗ����S
H������e��]%�ekS_7e�u݄��6bh��آ��8�@pOsq$���s�͛)q�_������������@�{@Ck!��b�"è�� O�X��=�ç� ��o�8s��:.�5Hc�*���:Y$mA��\wξX�}��u}g
6��v��v�ok�T�3������;�NJ����-��I+�*�ζ�O���]T/���h"a��9\�Z�,:T�]ܔC��d�KN��l�a�ɔ;�$���ehA��!�>\���uU�F^ڔfrAQ�� ^�k�񖳅8f�����z4s��u=G��!\as9���ǒ���ZbUl?�RYWD��N�G��l�����pR}�F���n�`��GȹpZ��B$����q�'}�Z/��i�;��$�HB�h����\�|�K�E�ѻ@����_F"��\V>���J�����d��N����;��c��%?	eNݚe�������������bHr�b��y�'<�<����CN������@@Wj�5�]��D�*���U�k^-Nn�A����-[Y���O�Z�����uS��wEF;a��c*�*�D��W;o���s�:GS��K�	�t��a������`�l��A ��}h��֚��D���;�$gYBU��H��ò<
�#h���wG�wye��З;ʀ��^y���)S�/�r�¶����`D��#+����q{�+��>n�ǘ�U&���u׌�r��n���`�"�"H�r8�鹎�!n`��,2�mb4)Jk�Ag�
�'�.ֈ�ȣ�4Y�:U�<�ucJ�3�cM�|��6:����42��i�t{��(���~ =����q��4���kl:3b���9��xG�9��|���^h4!��_�.�sg�g�b&/����7�O6Q}�?j�d�v^�T-�Z��e��l	^s�cu��F�:�ґ^H��*պ������&)-�D�)�kn�{) /v-���s0"/&�
�������z#I�Q�`B�7��V��쳄gy�B�;��f���D7
HE,�vl@9�^�j�RA�t�/\�)����E �2���n�ex��te�ȩS&�9?A5�]� �Y}��WO鰳o���<r6�:L��K{�>��
�^�3I��
W���a���Z�/֍��Y���d��R��+ؤ�#��&uW��J%�9�F7I8 nI;�h�G����<����i�j�m 1?�^��h-�IT�<6�K�9����K�0_�E��3���L������HM^٭�<���m�R���y,��Q���R��q�&�K4��pif�_6�*9��{P���P|��	~Wdc��>y�%�׬���-vc˃*W���[g%�� "��4j
h���%�c�8��ϳ̔VLW��"��NR8����{;��d��Ҿ_��RJy���f�"2���Lg�|m�nR��Ã�����e�����.�t`[�5�:8a�T%/P2��hI?�9��JAT�d�X�]'���/�폃��D���4ԍ����1=Ū$����V���_����p�0"��]S���vJ�~�ZA�F�La�ߝ���X�Eq�G�-�hM�u5>um�=4/���-�Ŵ������l?S�9z��B��@0�B�G���tp7!y ���ф9�]��#p(���z�����c��7\�0P8�>��Ȃt�nr���G�OO�C|�O%��c��2����N>��[V�
<�G�����@L&�$���K��u�`D2�N��y�8�ϓh��,v��iD�5��I�
�<�5Э&��ȋ�+Lcպ,Q��<�`�`cà���}�D�aj�T�(����r�
��9-�������)�}�p�FYj��e#�"�I�];����UԸ��:K>~p5OEo�Vg��Ý�ץ�͙0�
����7�"�Z���&3U�P#���u�]������߁�����񤰗D���~��P�4<�6.�Qb���-�6�rw��(���E��c�3�P7��"���Β5� ���e�����%8��ͨf�z�%�*�+?��AǾ�V��<]�����x�d㏸1>�|D�UD9��#42�V`٫��B�?)8#!��:!Z�w${F�1(|�Ve�Q\�Ԕ��u=��'gz(�a����X,%�砯C*W�o�����oM�	a�36*]E��ǁK��d�-�F�;��I�^WG�q�`���G���`V�K��c	!�Mi�2��:h'�(l�z�ټR�&�F�ɠVoH�� ŭ�F`�AC��Mô4ޭdӛ�]q �H�(4k&�+Ǣ0z\?0h��]��8(PLs�s�J��?�
�y �8���.�� �o20�[�ցs��>5�]�PWr�>�� x��Q���k�lu'{d{������&� uU��+���,��_��m���p��J�d���v�-��@;&%\0�����a�c��V�azY�:c�%y���	h�@�k��YL>��79��/��b�֩�{���1
�Y�֚�_Rt�M/q����§�� �uh�⹝^�S���$�`qH�)��I:vG��-͘�'g������� ���s��S�}�(z����K��%2X��{m>��-�F�/��}����j�Ow�+K�/n�������3T�1����JI��8:ɍ�׫2�S���Ɔai��T���5�O��o�]�V�vޥ�yzk�sZ�J���P��6�.�3�dd��{j�f5��.>���&oO�G�9i�>�ڢ%&��,�9�'�*��5d��P�5ËC��ұ���nbEЌ��
�����CJ	W�e���~��S�T��d��"~0���j��a��4����}aב��G�<�g{6(3�b-�fC!
|�Zq���O�|{��h����!��xk����d��W,}	_�\�M�àbX�e$��~��!����؟[�a���Q�Dɼ��1�IX1ȃ�L7'�����ނ�7"�[tZ�#8��-��`�률�`E���j�`ږЬ�Ʋ�%�GHVm��6S��7� �7z���Z*mF����<�{'��<��K�D�qLJ��B��0]A��*�uYͣ�Vs�&�����/�CR��:���f(1ǆ� ����W�*�#��nrҪ^�"Ȍ�����hU���]G>����Оn�PլnGxb*'��ɬ7��F�]'Tb��?���� ���'��f�2����2I�Sj��O�e<��{	�@u_[zL��O����`sw�Dv�~�^�K9��K���P��0�A`��BQ{��	�C-գ$�i���O�t<&��RԎf!�`/yfV׃2����xWH�5xǠ�<^� ��������\�|P؅*Ƴ���V����;@K�|����CQ�~G9[�O�8�C�rF�w^�(�9ё�U���X�̚���ús�S9FYR��L����wr����X}~V$c6PL&<Ց읛[=$��ޡV� "�xT2
�IMH()9~�*uԛĊ<*����š�'@�A֭��y�L��}���G^pY��X��ᬭ�ȓ��3L��@�oUZ_N�{TU�$����[�a�ul�.e{�.yc�хy5��ƩL�^zd�}����c���ӌ�>ɴ<�qP�Y��?��p+���������װR�[���{����=��k
���TW͑�����������Z��� ��_eK$g�P
d���#�[C�ް�c>&�mx��i�S9V��lG�ƕ{d���9�jO���#V������@e�$���T�Z;��5�InE�ʅ��ja/Ш#�����yy���
(�l�
�|l�yG4%��c��xu�Y^���s�(,��];#�������<��z2�!���@-J��	O�j����T���聣v i(�v�4���P��v��J����ȇ�#=Ɵ���ģ}��m�|)��L����M�)�� nP��n-�e1~�ʑ_���V4��C��wQ,��{l��='�oG��]�X�X��e�F }��r��W�"���Iҙ�F{�լp�Н���V�b�_�^j�4�W!��fZޘ	jc8�vϩ��E�uҭ�3�g�[t�G��/��\���W�	9�ܺ�Iq�u2X��拦�(3@�f(�y�����E�-$�*n�n ��d�f�
\�˗����vȤ�P�n�MP�����6�d�%?�[ZB^w1ߋޫ��S�6е���ﲭ�w!���x���"�hJur�R�S?�Ov��,� h����Ǉ5r%ʼ�_u~	�SI�͢y~/�8tV�l^Ƈ�i1��B�G!kl��<-��|e�_�����t��Z�^�����A�*�-��j�K<��U�#����é6?�U���B�5f��E��A���|i��K������[
#>y=Z�('�3.��l� �:���JM�	+�}��]�C��'�2}���]2��5ͮnXw
%��U�� �ʮ���g�|��v��qr�
+�x�u�l�ѱ��?�8��&����[V[��a��-B�e)x�ȳ4_fu����%����ַ/`�N/+��ip�X��C���R���`�Ҷ�&HD8&{��W^8H�n��Υ?��+��F僇�p]�Y����񑻂?�	��`�$P����w�yor���9�F�x�UO�WZFs�T�����#B�t���UDt��C�o��#�7�E�{�*�~��z��8",��ra�>z{aL�$ױn%�k��Q�����:' <(�͒���jL�p��A��ȗS�q��CE�ƈ�w������jͦ�P������4��Ϧ"��	�5�0�*\y9��n�_.,_�٢'+�pVzl_�/_`���ܼ��S�(ԹH����x�R��e�`h�,�S���Ɉ�����<�z����߫���7~{�S62�z�j�$�y�;�����s�9���-�P&��V����~��U�4P��tA��FxqQZ��:�1�87,����L/૴�?nڅ����n�L4��Pz<Nq����X�,5<�ǈ�n���f��Bt�	��(9�
��i,&u�ǓR��4.{���+^��"!��m�}+�kW�1�����~OP�)/D�,G��xwW���E�Z���Ƀ���<���.�D��˃�"��[ԟ�M������&n�v�8�0!�Y�����pb����^���z�dY�l�xOC�>5d�ƨ������^C��
�y�����:
5�)��3L�E�z�A��Q�������@bx\�/�T�/���(��ܩ � ɏAv�6��&CP"M�cK.����=�YZ4c��i��d�8��b�O�ЃBmOkgD�����q�k}����z���sd�dE��7��W����ۏ:����t�Y\UǓ�c��2k�˫ق�������k�	x�o�ߑ:C�g�-�����G������vBm�Hî-��!�褕^��h����8�v �������d�WV�����?�q�����(�pa��)�"���cm7Kp,}�B��-���.�5���vu���ݻ�Ĳ��!�׹$��[|�[׮���<�4l��ډ6��g��P5�(�Q��t��j�Q6�
p6�(pQ����/���Q�X��`�΢��eC���f� ��2XN���6+���#@'΅ws��~�1C�c�f�Y4*�����aJ�����ɞ�2φ��6�#��N�$<SΔ��ԗ˲���b:S��r��4�W3!i��)���q����:����M&��m�h�������dk�����zBf��|�޼�l�̆���\��k�9>��=��!��SA���L_Z(4N�#)n3�yX(�Z!Z���[Lg��?�K�e=�]�TnF��Sil��S�������k��DEkӅ�~�[�����?�
Ɲc�t�0z"3F��g�q�6~V	�#�����vO���J(>[�<��'o32�O�J�
*� K1@9��9z�2'`�ӿadh8i�a�@��5$r�,��`x�C�(��Y[F��yu�'�
�v��/�$�Z�m�����?P��u��ȁ5�~zʂ��W�5阀p�v7�&�m�ۂ��0��o�Z���%d�'��|/�/Κ��ٕ�<3�����B?��W8F	��&��E@��� 4;zҦ�H!��Ur� �Ŗ�.+�������,0^����S7&��w��}�.w��g�o�.����ݝ;3y~�fC{��������)2���)��Y���x���:�/= a�+���/�+"�a�ÅV(��K���J�+��HX���2l�	C(I!gtz��:z�a���Y��0��/.��=�Ӑ�T���g^���x�4e���+�z?+��}v��eAzB|�����H�
�)^B�O�g%ŚM���~��j�~Sj��?�Q������]5C<ӡZ'�^��+�<q�(�u��]�nFC<�s���»a�`^��0��n��c[�����N����_��h��P{(t������vC��݊W�r�p����zT�;G)c��{��J�U��P[Q=ТA��,+3	u/q]Ƅ�2��=�W@�� ���ǎ�q�?�O�� �|�1`�&�ޮ<Z�ǗS��X���ŧCBC��]�	{)U"�7�^M<��r+�Ԙ������e����_g9Duu�U����c�G��	�V����6��B��?p���R�����0`�.���eV1G�L:��YwZi��̜���$�8ںo�����W(�Q(*"��3<V����D���^�)h-3�E�KO �a	@ĿҔ��:<��a���/�@�uK'X�3�&��,�[�n�E_ ?W����r�X�&��������/��)4��{8w�<cև���h8��x������'�9����C$�����b�"^��נfyQI����O���E��ď����p}�LN�<�����u�`I�g �<���$8�����!�LQʯ 4�4�zh��bX�Y�+Ċ9����
6����$��/�@��:E���6��J.	\���:��_����e]��?T�##�I�c)�B�*�#p�ZObք��-D=��ɛI\���L	�l�k�F�<��j��ՠz�H֡�M׍i�V���6�r�>�n�cȈ*���IE�%i�范���夾��%抔5��ʹ��}�H��;D
��(ϋn~��q��Lg�"�xcP`W�Õ[���Ed� ���Pi�O@pA�*>�S�d<s0M�`Bl���I�i�ŗK֘bűůx[�!P�͍?��E1:U�vJ��7t^^���������=Tй�G���O�K�,t5��_PF�|pN�u��Z���u�x�y��S-�Ny"�8���C��R�*} I\�K��-8�-�Tdm����5�d���0�U�__�u�4Y@�E�m�É�������u:�y�1͓C�?��Y#`8P
�D�0!��D��`��@^N<�%��7��ףu�C`�J|? ��!'��:t�ԆX�:W��t*��'�H�Q����F��vҕ�~���=�pϠa��`PT���Ы,jH7}K'n���Y�ZV��4w��|��m �tK�ՙd|�$��^��	�鶓�6�x��C�΅�ʻ�(`����u'��I�����l�zTDA�����0o5O��L�����	��0� |sP={�`�\`
3q���Ԡ��h���d<��������oU���^ m���*5?w���S��f�����#qF���ac�Hjf>>]��QH!�9S,�����M������JB�[��Ω%��j7�b� � �4�����h��v�}�\(�"׵OA(����s������ks
�$ �޳3"0E�v+2�����˲h���N��6� ���ś|��	.��I�8�y�[��=G����luf�H���
{Z�b��
, *��~9���x�|0�����"�Y�iv�.FY�ӳW����NI�Yv�T�DHNՀRپ�N��2�"�T0�]T�27�{��'/�]o���.󄅐�����7"�����ҹ��³�2��Ѝ?|a2i%§Kۏm�%�d#z��i�=�_ze�K���FJM�b�ny���t{J��M��Y���S£�!�6X��a.1��0� �~φ�Q�$���0X��z��T�~Lf�r}Y���뇨`�&vX�e25�6g#oC�S�5���"RT�	P��a�"%��^��¢�I0�,C�ٵA����_1�r�加��+w&~0��v���gC)�%�ܣ9wxU�-3xHVV�q�.ki�B���M$�B�#�ۈ�ؚLǨ@�C��,$��HK���"��4e\E�1�)�sׂ����-ܱx��Y�=]��Ӳ�Mݣl��ۂȕ��ܢ�j�垞8�y���C���dNB:e���s����Gy�X.���Nfw����<E|�Ja�ͻJ}tOC������w�EJdѳ)Y�U �e��PJc��A�2���"k�߫�^X�+��*p������i]���>��B�Tsx��q��/x=���E 4�H���xy�k�Hi�y� �.�(�]������O���^��PMPTP�fBDte:ɚ~ K�J^�ovԮ{	����[��Juu[��o�ca�
�^�V�u�0��*�Ի[ܵK��3���K��u�F<r�U���d�|��i�G^)��R�Ȑ��H����V嫇�L.�i�סa�P����shECޗ��Ϫ����g���^�j��|�"��[���F�'��(�b��ݭ�*c��y��ZP��&�-~+u9��zp���0]\"��Bf��E3��pt 톆j���Y����v|�T'i���=�&�s�77��oZ��-w� �t�nI�t��*R+xm���D���Z*Q�� �<|d�4���PJ��W��L���r��A_�U�e�#�=�j���AO�jfj��W~�j�a�S⤫� �LX2f���.����ad�X8Eg"�t���Q{�8�q䆠�3��m�����w�-�
�Ԥ]�RS_o�!\梃<���\�ýc�y$�U�l4C��; (�#�2�`[�q�3�٣3ݤ �mQrV_Z��x'�(�t�7/r]q2�4��{�^�#�9/¶� �/9��Ԗc4��*p�.!�";lM�E%>����R=+|!<�u��1˗��bG�!�!9�ކx���r��F���]�U����]��E��0�v�MG�+�����z	�N�z�u�<Q�m����cV�G_ҡr��C
<�;�2S�8!��}�\.�1D�����_|����j����`n$� �����8�ov�y�(0���8��4d��v����|T荴��ګl&�г�R�c�:O��m�kx��i36/˽�u�[�|1B�����}�#_yl ��� �	,#V}yVi~�{׬��C�f�]�L����	��!��'���x�=��`��nJD4�^=�<�t��ޱ���ޗ�a�>� ��La9�V�˖xR8�XA??�:yq
��N#�$vc�����$����ϋ�41`$]>d���d�?����ȹ�m�#���+I,���6	�J�T�'!م����&�Ϭ��v[���]�'ST�[����p�<���2� Ain!j��g���I�>�Y���i�QB�nv:nqM1B��#\^����%8}B����6qQB����Ǭl���c�[��Qͪ�6?�>fz��'bM�͕�!��>�k%���ͩ��p��v����_3�s7�"������G<�sĮӢ#%�x�H��T�Sҋ<���T�k5���(�����E���9Fd���rG-�s6TC^��*H���T��͒KM��ӛfе�{��\ eQ�D́D�B���eB�$-�y��R
��-�'S'��C��҄��݆M����J;J
�v5� �~:�R��� a#���:��&�1]@<�R6E�@D������(���8�O(�z���^�G����뿯����¢NXzu?���D��yT��5ˤJt��	`H��s� `�> xE�x!/�,X�I����/�s����\��"������kR9;�K&���1@)4�fs�Z#D@@������u��h������wV�؟Ɇ���N����:V5�-�|�lmR��� ��艈e8!���%)�X#�a�L\�M���;@R�&4Zw]�ĳ��K5?�F�jH��7<�^��M[1[����r��~�v��'�R��)�7�� ����VFӔQ��)�zv�����3���p�S�c����'���&�_�ѪL���D.�*�e�oB[vSv� �����F�B�a��F��E`!</�`�T��k�N�əh��-�ܰoS�����xN9ω�g��^� � ��`1S��|�Ћ����)�"�j��ן�B+�t�e���Z�;b֓ |_" ���Qt���_� 9ڔ���:�i5��<a�����g2�#��`Ï�4_7���w��?�S�3(@+7��c����l;yW���@��=��Ց	�s��h*o�74
G�F|Vq���a�*͘v���`w�J;��$��5]W�A��)������`�R�.��~�G�Bb��Y;��l�XH�Z2"������hY|�HV��i?����Mk�Ѕ�ے��ʹ3�)�8F�8�_'�)&|��Ϩ��|��0��~��u*��s+�'���s�CC���
<1��1ն��J@U���y�@�J�[*����f"Tqm>���>�{:��B�f���,@_z����E Gu�^:w@�_m<��]J�y��UD��kff[��l�x=�������mXҧ[�)��qYڵ0?Ym�ҾK���G���Z�+�^u-{��֟��ĵ-l�
�^Y�]�[2���q�GL��qU�Ͼ�29�I����D!�͂B?��_�_D�^�M3�B�p���О����n�՟�s��O6nz��jS4�`*���lQ��#
���Z��:Ƈp�ӻ�+}�r�/M0�N-����>��!�ݾx��}Q	�ۉV��W�k�t�Dө���zR�?�\V��z`���T�� ��V��� -�z��,	���6��=��qb���C~cS ���O��l��
!�����H��	���A�n��߷�U߫p�ȸ��h.��f�K�]s:����:��Y��ޝ7�������tk�$�i9'�J�7��Q�Hb���>�<���"���*�ݠ��}���p6��D�Fl��$�l��Zy~V�L�ڬip��W��V��:7�tx �>yP�L�7H�q|�ˇ�L�j��Կn���ʵG��d��D�mP@�d�lN>�f�$��س��|�-A����5|���>[