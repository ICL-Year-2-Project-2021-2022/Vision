��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�@�w�4�R*��D��*�j�ޒT��G<X,���4+����P��at�lsR�����sm a��W-�e%xYM�JX�t�yˮ���m5Ī����;�"L�#R�݇��y�7���i/�5z� 3������a�U�G�=�mn�Q1��wԏ�%j���;}f/&Ǡx7|�=��s��Fܜ=�y�f�w'�O��g�T8��JIV�S0��d:��ʐ $��z�,�Hָ��Q����C?�J�0
ֺ;��tk���g��O���E�х-�e�,^���lӞ$�Xg�p/~��+�o�4A��޻Vȧλ�
ԝ9}�}}[����/��g;-?�	�kF}�t�~c/�F��<-dX4ƻ-%h���`3:�Q�p�tj���6\�����U��".y�Ss@4�~{��N���k4�$�)���F���P����ZƱ�i+]�ҥ���-EđT-�qe���(�2h��q�f�f`ո��h�� ���
��|���٭����o���:D@[Р�������x$~2�j\'�n�h��^*j�fH�.�&��ϣ;�E׿���J2���$47GT����d�q���mx')����T������@��T-��!��ӟ���`%{	�B��ǫq]�K����2C5�m��_��MSr���d�'�0�^-�o_tvYD���������o1�wj�F�u��mƎ��e>=KC}'�r%Pfs��1��a�wD-)v�/�1m���pʩ�=�0���c���RW���*I�@�a�Uޭ�V}#"�a8D�6=�p��v�@�K,����̏Q�=:zL�����u�򓁗Z�>l�,/������R;���SL}&}��u�X��EZ(�Ӊ �;߷�����C��L	� v�7��k�,�C���PH$i*�Ы:��4Fp�:�ܟ���.k�>��ʟ
���Z��̅7�<R��l�9�dVX�f{
�t��Q�D�ͨ8����Q��_��oό��Ukb����Z��8� ��s2=����Vdv��6o��GJ�f'M�æ�����n��9����:���s���ۛQ����sS�>Z`�q�pT��z�'���;�178MU��>�9jK�q"G�v�x��ʹM���.S�m�"���:��8?ױ	��u$~�W���h鎀T�L �vչ��R�i���Zl|w�%b�Kr�У�=���3H�-{MrZ��C��1@�����(W^�8EY'�=�'lU�{���K���.���cߥT�����.�@��SbgU4D���&�u���z��%���g�Ƶ!�E��|W;��d@��a�!K�V��u�BT0�;m�	r8���1u&�5��f�T'�g  #�A�'���c���ғN���P�rt�}��N2�r�|�:KG�����H�����D��DJ�����n����X�2�,Y��I���Fi`��s#�FV�MM�}���W�r5j��֔ϘB��ѕ��Hֈ�A��&rb�8��@ɹʰYk���v9zT��bQ��52q��B4ޤ�׆�!=0T�j	S^���7����w/³�w1�*�2�H�׬�o�������35�������h�G �E�
���e֤J���Տ��0ѝ��Z� �K��ZmN�B��� �	�W�t�������;t7AE���~QJ�<v=W���R�S%�-l�ic�\�ӌ�B��Hu�N1o�N��>�|(ddfr-��^�>���y�q��V*��F�����Ծ�E��N�z�xV%W>97}XX�H�� ��g����]���G�S�����5�5��e�ZwL���lJһ,g��q����WR���ߌd���ڐ��Ti;��.��#$T
p��?�K��B�g^�/�⹥t�eG%�N�C�0 �Պ��n�_�X��*][�c_F�,aQ��S��`N ��S�j�ݟ�v�̭���'d����X$nh�S�X���O���^rL=s��n�7p#P�O��s�݁Xх.	Y܏���Q���Nu�q��6y��=]�u�8k��6���r't<�!�F���r��"���1�y���p���I��q� ׳�$ͳ����!O83e�^u���+C�i�Z�0�Fsg�!�2૯��
�ߜ'�T�8Tq�u�^["��Fc��$�&\:hp�v.W8�r�7�\�H(e��l��=��N�X��a`�F��TS�L��T�/�a
��Xߺ���a��O� p����qA�hb��f��P�rYO'�^'���bAb/l�:S�uj�%��|S�X!��q�
 a�P���.G�ª����>&Z ���i������+CR��o�����Ʒ��)G��r���U֫  �sM,��vT���0Ȓ��A`F�bF)�eAZzx������ٻ��;]��C�N����5t�z�����
����PԆr����U
�L����k`��yyf$`B�F��F�7m�:�z��<���C<o�;�[��<#��<'PRa3��n������!�D����6}��9�IX%���V���ޒ��c�2�u���!��|4���P�W)��U��,e�[xcA��^v�q�#��E<��p��%~�5'���o��0��J�F�.U�x�3��m��ŋ�%���4M��W�O�b�j��<�;tPPu��"g�TK�2.Jܖ��k��Ri��e��7t��5e�����>�JD)h(�\�!܍&�����,
��{���-!�9pf��%���7O���9��V����ݦ��$3��B�=�
���-`;�*���"0v�jh#ފ�a��-Sa��e�X ����=I��f#էl��k����B�/UCW8�Ƕ�.��:�l��O�\�o(�:hn��7~�FX}3 �I	)x4rY�v�Q�C�5��z����G�4xd��w�G�7��LCΥ�hώ��c��:M^�!��^ny�<ȴ0�he͆H5Q�[�|	Ƣ�jG�w!�t{�Ȯ��wݽ�pns��C+NY�,��4h����K�MK�L�R##�B�"��x�_b��� n�4�*#f�����%�E��b?:�H�x2�s�`��C�����aQ�t"��/���+o�s�J�r*Z����L�Ϳ����Q���8��wi�c�P�A����*��גxI��{@��Tg,2�1݃��V;��$�.Z�uܚ�E��]�&��t�$��L8� 4��Wr�T�[�(�~�o
^�d��]�A#{(�X:$Z����~{���g�K��&yXֶS!;㍯bv��L3x�|�],�a�큤g���@q�����9���Q���N��13�¢M�&�V
}��k�l�^�'FtЬ�a��Orod�X�U�f(U�ݠOK�|��.(�1^~2b�6�7z�L�\��4���nI���u��pNԉ���I�<��D9<%���#�
6�(#�Y��b!����,_��;��E���pvɮ��P����(�W����n���6���n��m`�VD���
�QI��@�VŘ�,�u�3'[�ѹ��=%��"��M�`�����ڲ�R�2��$��[�Hw�'_���+`:>��<8��3����Hv��\�C�e�4:��KRrii��Wu���F�&%�C{��^<J��Ȝ�1��An��4ێ���+�(Ux��&�M�$T<���؈�	�Y1g +��������n���yA(>�j�pf�����֢�. �S_;Do���`��fF��&y�b����(��Q�v\��f�1L�p2����뺺C�(���������U*v��qg�PK�$��΂��_|��I`�Sr��өb�����"�J����;<��6+���~�S�X�^���0!S���o�3"e{)0e_�&[LT���br`��	�ؠ^ƪݮ�^�hkzmD	^�'�ȣ�����x�� =<)�m	���)��m����J��� 0��DpŪ;I��cդZq�i����h�L��Y%��_���y�nh�M�Ջ���	tʾy�v�}���t�?p>��g�ԡ��_��{�����}�IN2����
1�WÌ��f>���E�J�l_�`��>��|Ga4�N��%�&z�=��$RG˚��Wd���!g׎HR�P8 R<B9�6�
6���1���b��ց2���� �/Q\���Ok�1EYq�s/�����߻�f?� � .��ӽ�x*���5��I@���l��N2����ZW��5�6�;���~��V�N��չ~��u�G�}E��=�8� (��k�f�(��o:�W�O��An4�8<�au�gN�-�#I��k�[}ו�!ŵ�>�yF=?�m����gQ��|�<��ctɳ{'�q�g4N
��u q,[���Ԛ�,����Ei��X���X#�����D8�8��������K�M:]V�=$���)1m]�&���ʐW;�5n"�g���y�SW�~�>�-��SO*ذ���Mɲ1s�����P��0�B3����t�S'J+T����>K��sO� ��Y�5|��u���gdx��H��Z����X�6j?�>9~rN턓���b_��X����,�����6d��"hV+�I�J��q��羪��9���y��-\��'Ԩ�@�YI*�Ɵ��]�T�3T���̌��8��2���y'M �@�;�I��:?��ڳ�f��K`��{�Ƌ9�Y�� [0e����ҽ�l�ri�{�ʦ$@9� ���%D�4!O���}��v�-�X ����2��R.W�VT3��!���S��	��_H/S����n�̢��-��y%�����0�S(�Y�5�Y,������k=���ѡ�p2�.��tn��CW\h�F�r�*��}Ц�l����y#�عH��}s�|!�U���U08.Ѽ�	+æ
4��юyb����k[���Ze[�|���A]�%~��U���\��8����&ލ?�>������t+�@��{���{I�qi��,/�R�?����ao��k# vHO""���x�T�*q�5�C�j�Α@��=�p����'_�-h��)K
D�
W����7�v$d��<��4�q0�^�A������
��$�VU�a&��8�~&b��cV���EI��qF0*��ī<c=�^�������*V̔��y����X��B^��Qn���p��E�����u(Y�Gl���ߢL�V4 �Z�*oe�����譝6��d�����b����e7-[�;1å� I<(�����ު�2ƆQ	c
%�O�rFZÈR�MM�0qG�ܲy��
E۬�o��.Fx�%Zm�0��HBkA���B�t�
�j��ճ ����Gw�<����Ź�l+���f��PJ���V>��hzd�Z�D��{0�$*����8��7p�o��Ͼی����6�u��8�@�=�/�DXj`���+����kKt��0�X^�;��ANW+޻j��{�ExVi`��/�5��A�< zI5Z����UD��O���6@�u���R�ADM�>?2�N����~��tᬧ#�g��jn��`B�Z�{�#��#O��Xb�ol�,Be�B+X^d9�MZx�� �u/P�jT�|���XYu��/,���Y�;.��cX��ς�X�3�� (��쨷p�GY��ٟ
ƿN��b�:m��Z7���\��| ۞�(� ��ԩ���i}Ԓc�ȯ#,g�ID|-�NęT��sI�1GP�C1ӀQ�x$��m�EW�<rl����� �4�p��Q�C����g�)�R|����7(���C��+�)}d/8u�~E��2�a��F\Edv��F�ӯܔ�l�J�BW��eÌ�a�����g��V���!�@ݏ�5I{�w$���H�1⡛-�0P�O-{���`�%w�߽ �[~�hя���~��� ��x�SV��S��}�N���H ������d-�G�ᦎ��m�|Se�����*������ϱ߿ۍL~l5�6z�щ+���F�m�l/�G3
;C'��:��UI�ne��=�M	Y�cp���m���޼B�g���[Uy}�0�h�X�ng�<N�����
��Gn~T�Cj��%Oh�Y��qA;G�o�v3�!�EEf�Lj�,�αW�k��ה>-z}��8�\�Dx�d6w��/y��*�K��q�� �e,���U;M>�������}V&�!k`�/6�l�������Z��i7�3�˝G�o����iA9�:X�U��Gޮ��)�.��?�`S��n�Ƽ�u$~!
�S r�D����h�-ajbO�Xz (�I�g�W��� <�ߏ	W�v��W���������IJ�-�x�'-:��T�X�A���_���Nv�qw)|�
R:�8`�ݐ�)ﵥ��c*����
���ʎ�z��ײi�M��\4���=��F��*p��sʳ�<��&����W�5w��n �}3��I*����x�1�Sּ,��i��:�(�]�?�{��9^k�f�:�!�}�\sZ�`�d[\$d�9��͒�w�R",y����%!oD�W��Y��T�7�t�i}Ud��WE5���l�e27T��rAB��H`��f.E�B��Z�$1�t8n�����A��mkv��0,�+i1�A�}���_�#k�hw(��ݫV�t�Q�� �_%z��PK�^�4� ��"hz�|/"6�2c+Ismכ��f�X+/��Du)���@~!�:��"����Q��O>�w��CFj���x��l��O���3��D��G�>�`��ۂ�w {r�|תx�+d�%��J�����C=�펏��&sV;��B[��ڔa�xd��&�0r�ܥ����a�~F��{O�0����S�pEg6�2~c�Żg�����pYi�ɩ�ǎ�;18����T�K��w���Q�c��p,D_�:Ͱ�����D-�@+�ˢM4�����6�8+�|��>�f%�6�kW��)|�PO����g�V9<*k�[�����mn�4%B�h�+~LL��Ň<�'��h&4d�0�����<�k�[�%"�P���'�	���%���RoC.lV��l���(�@FZ�^���J��Se?e�!�+Z�i"����4|�M�1�=P����D1�2�B�hL��Z�T��:��n�9����A��ݐJ>�t�o7Cep� �}1�aÆ� �~�}3��M���C?��6��;��rø�Г�E����i*��m�J�[�+����-=�[��n�`�o�S�ݮ��]�^ȯr���6����D�:�I0~"���䭰�s����<�G�1��^�{�?}"O0|�X}բK?���w��t��.?M�_����S�W4�Rf�-��e�53��k�#�Gǂ�Eږ\Wz�vF{�mz�$�_�m�dD8i��S1���rwB�Ǯ.ym����U)`H;�uu	��Ƀ��KN�so�nL�?,���A�
!��m�}�tF;T�r�����ivZܻ�Ҽ��6�&v);$��g;�mt^��]P�7H�K�:���0��F�`sC���S�+c8C��\Ⱦo\ �����]�{�-��DI�������ѹ���KN}d`�S%�l���aL1B��]=�8���lE���"SQ�F����?��eI�/�b��N�C�.M��¥����G�Ȫ��8k��4��c$��N,_E���??�?G��?�=��,�wq���π���s��o�z� |�9A�e"HS��s-Y���utSP䦋�3k ��
�r�X�����Ye���~���.4�`Cv���6}̈́�s?����G�K:ic�
�v���X�D}�Nf|W��^V�s�a�Mñ�_���×��ycѬ�Sn��{�$�:M�x�;%9����dV���p"FĊk̫[�t��������,!�)݇�n�癜tD�C�m6>p���
#1��H�}�F�0(���F�Nz�
�;Q�5�HY�!�0�P�'��d~�j�L²M�WIy�:F�H��� �5L~��0������b3t[�B-��e Ř��MV�w��$r�.��]�A�,1`<[M�W>�2-���f�Z�?Iu@����7q�r���FQN:��6\x��ht�6�ˆ�.:�r�b5zm=���2�>Щ62��ܮ3LE��$H>0�!:<v�aՑ�}��g2#�'�/,g:|�%��&�52�st�ZF�߬3��S�b���v�W�0���U�a��m����-��$���p*�T^�O�h�k��9����//P�zj�u�>r-br�Hn�KW	��@²U5eν��	T�-�;��g������x�=}x��n$�q��]z.�]<� k�G��+fj��m����ˊ�	�B���	�N,�)#�1����N���*��g<�eH`�n�$lhG��h�.��u�V}g��W6�XX�GKD���`����9a^�r.J�xc氳���HRtW�QL_��y<)�+��pa��{��Ȉ+l�l+PKj� �H��֌zyO�xӪ��}�42Oʰ�Prp~ː���r�>pm��-C#�>q��.��=������r�P�<&� d�x�]`(�91���/�RեuH�c���J'�YI�8=�p2t����G*C9�ʢ���9�,����hoP�<��N}{�j�u{V�bjY�f' �R�mƏ����J�WG�Y:;E��Wbyx��q���E@$�*\.�'$��<�AZ*$z!w.ÖB��٦eێn�o%�伏<}���ьX����=p�:U;��Y��Q"�[�#~i賹��o���ք�ͺaC#R�k2�a
.t�F�Y��N�e(�"�����=�v��@�o��O����k��N[-���́ϣL��6���+�!u��7��;�ߴ�o��v��&��:��4��֜���~կ���ݚ��b�(��2,1�ص%�rC��)ɻ�Iy�S��#�w�f�w_h�
�xz)*��o�ئ���`@�)�^|��5�J9�������'
���`���f]�K�f�4��c�oB����z_�,�lb��+[��%dN0�i�v(b�?�
��eܑ�('��\��N-N��oW���e��?��*���9�����n��#�B�d���I��ҧ7yN�q՘NX�z$ׅ�������[�:��ZE��/T� +)��C-��#�[n蕑r~҄���taޜ�}�W�F��L��8(��-fk��$�)&�3Tv�&���9���(��lH
B��l&L&���&��7>`o'���ɌC�OM��S����N���;�}�8g���ؿ>���d��:Zy���#����K���]��GO!��l�qa$�\\�t?��/�:!����z	�B����?k�?R�/쒨�ǵw���.�C��%��(���o�����`#�SJ�� �����߃����Ee5�؇��g�şG�-����L����R�~�d
nEx#���A�ɣ�Aۧ <>Z�z ��b^ñ��
����J���9,A#�$��f8|�0�^\=\�qYIW��B�;���A���67$��M�x,s/�)�:U����l\{��Q��U���{	��E�; �_�0��Bu�o�:�I�t��������1�X�X�@���0х��^��p"�N����w�O\Mam�Լ��2�ʺ��[�q�=�}��"a]���ZN�Y]��}�-	t=�ǒmM$�t:J{�����*>��ؚ�;�x_��X���l=�4�̹#v��a��r�Cf[���G��u="��1��Vg�Z?���Q���k�D���7�����o����nG1Ti�7��	6�A��R$b	����6c�W�-(��)r�YJ�@X⵷�YN���l���װ�E��fja��+���BĤm�r��5�esּ:����з�h]_VH�}����ll3Ԥ���&����.T%������	Y���[�3��F|������Ff2�� <{�M��7���-8`��S�̀H|�
O���-LeJ�qdw�4�Z�^�ES�����jzIou�e��k+
o�K�E���ݫ�S��;<(;��V��Mz�7�r��*�ֶ��
Q6ߚ��%5@������aX�	G2��D�������u�'h�C����l��xdDyh��U�&�FPn�ʶ��d���W�R��_Bk� Z�xW�����O�9�<�C�ojO�b�Tԇ��n�ooD�/S���bY�9�Pڴ)x�R��#��x�}��Fg"���B���B��nm�DpHɄ�U�rdwN_VJm/S僮��,H��X��X=MV�s���?d���Phb��q�N�x)�ж	_E'���f�^���N���W_&�o%+5�>J<W��v`�q;��n�*q���lA�J8'Q�1���'�k$�!4�������5<�>e��;2�d�=m�@�:�<]MJV������eiE<�E��������n5R���p͌��~tI |���I~�8����tI�z܆ۙ� ����p��kܕ�7�v0���
�����^'�Z�R`ֿT��K㙀�-?�1i�Ԭ�n��3~_�^�j�]���]Ď�J�ݻ�dβ���9����k1C�����=���3�t͡��교��g~��*[e�Z���Z/���L%��#�yvz��w9�k��O�؟tY�0_g��ܒ��w�$��6c������?��B`�P��╺�L[M%���}��"nr��ΙA�<w�}aO��r}s]Tw����sX���`���1ްĢU]U����Y<�v� �u��OB�aA��ؠ�T�	�ǧ�x6)�p�P��ڕ9�X"���vg&�D@�{c9�k�����:���Q��<��ҫ�N�����o���o�C̝Y��Od:C�r!�[�E���`{'
�(��l�q�5��ԐK�;�&�ip�8'��E/�ʶA,@����0*�ާ�9�hu*���̅�y��i,��Z`�u�V��@fHl	�r`���qr~��PH�&� )��3+�6@�y;��������
�z=�Y���~gɏ���|�D�c2��^o��	��]�s������>7-S�x�C��V(?�dc#,D���
�������,�Z����0��D��uڳ��	E�+��
�<0�ۚ�7n��#.�ѹ4Bd���e�*^��W��^�$R+��������<Hb.��*����8���_l~��ʌ����a|P���ˌz{�VLN���5IA.�Rȗ\N�1|�\�fu��pU�0z�J�tp�uR����^n3��Sj��8fϿ(���˖�f���M�OӨ�n����s�����gq�G؀�A��m���J��^�a�d�+g ��g^P2D�zF��[��8:�dz3CS��@U*�O���Uㆪ�����ؗޜ-U{ �?TsjE.�ܓ� %yT*���
�(Ne<�W��h������qR�vxah2����UAb�LQ�
�G�n�>�����2D�����X���`��x/�ۃi����5��j.� �:���ӈ(��RD&������7>�yя$UF}=����ܦPFF1��J�v���P��̥���\����xj�+*cmUn����|�Q<Z]�Ka�݂)<����R�I������������0*+�p�4�0_�1���Sg��ʠ�'Ë��
�:E��_ǧ�)��4���z�Cۭ
�h�=#f�n!�Y<�io������c$0(���AQ�e��>� �}�W3��uX_}6P'w����*-T\��\�3�S��"�vi��r��B��Df؞�8�>�CB����渎��g#�]S�@����a �걾XH����§v��t��JO������@�+d9�O|x�xڮ��!`����F�+S���1�� ��^.�e��dm�nXX�vo2"��m[A��kC�4���Pv�r(R4���]#�֘� y�{OXZ-�fM�,�,�{������S�4��{��(������Sڐ#��t:� (m��/��<Ծ�;Nޛ�V+k���n�3ϓ���L��k� ��u^4�Z����%zcP�_�˦��@�[��
�ߡ$d�钣�U��I�����v핣5/J���ŲX�+"0������Gmji� 5�T��M���q߻nu��oOޤ �C�y���GT��57BךT[Y��ަZm�@F� ������/ZG��u+�[ËW�w� ns\��8>�Id�êuF����.P?��9����	j���=�t����~qBa�3���//��;�w�X���xė�(�*��8a���C�4�(�,�
��M��TQ>�:�bD/���;����@|�B��؋z�ѿP�;cJ�#Zl��w�F���Gj��9���4�ǘ}B�����dD/$b��)<�y" ��vD�����{[�����|�<cBȲ�����Q��c}N��*��\7=~&���A�������A�-B/a��K�[y�|�z�S���-�|b>�qj�-E�;���%{�˜)r� ��PR��AJ��ָ{ǢМ����B��z��,x'>��A0�W�[����]~<��u/n+ٕ�>F�P��3��=����;�߾��{C�R}톼��Jc�+R�{�WJOܢGWm<{EM�I���O*�J���[4CuD(�I�~(�C׻E �8ꜻ!֊�����ae��n�R���(�&�����!fg�^SH�a�[��B�<��sf��@�B���|�z���a�y<��z<}x�M�i��B�>ʣ7で������-�mSx�>�l��C�-7����G?�3��';4�'�I�9�'_�!7X�m��B�d�1q�+X���z������
�]؞�ǨV�e�A	^X�[l�՝�z/�ɽ�����O�B���C��q8$��ю���G��{���b�-�>2%j	��3��D5�#�Z魏���3>>WJ�aP������BS�����m����g���H¸�%��TyЗ��m_S�v�����\�{N�&�g�����7qo�5
�`��L�9��}��i�2+yA�Y��ݍ��<I
�R�q�eC���`^�xւYn�;	�9�����`:}�er}]�aB���,;��i�*����HT�o6�qR����VEѳ��@�)<X�6��k������܌X�m�'~��*����$Z�R��N��'$�[�������������'�Y˕AE1x���̓t6����m�=;=muJU�1�
��9�����q{�|eM��0g�$U�`\��u#w(���W{�������]��fE�t�^N��s�K�>���>��|�t�Ij�p /�)�mFV v�N!���}D���{>1�����&����i�|�^�o���εTH�X���ܠ`%D���+1���c�ʾ�ɜ�� IR�J�I��:���A���|Q-H<Ik����b+$�㓅T=�&)9d%�,���"K͙9֯�_���e� X#�Q+DP�ǎ�_P� m�&v��x^���W���&^I�z�����,hx�tG�ն=ӝ��;Ԁt�8��\z�zG��b�椥��-7j����/�D]G*S�d����TT9H�,�,7�X�ww1�y+���ȁ�k.��*Q}���h?H�p��y1�rT�l]��e�d���/hb�kp���9Wm�d�Tm���tE�K,�� �J�h3�����B螥�n_9[&xe�Oz}*O�hD0%o��.N��B�d�!�Cu1��C֓f<�:��u��|�ї�4E���G�?�̃��}�m����R�ݾ�R􂫵�nK�tm}��A�L�e�`4���|�ط4+��=�^�'fY�@D�+��屭Px���{G��m�KT�FN}�Cn��:��
���4���v�jl�.�����&��my��jeo+"�>�¤�ۥ��^�A���\C3��Jg�ɧR�~���=o3�"|t�/�'g��겗��Z8%W��� ��:���X�8ᲅ�^r?Y��u�.��*g7#���8�+���
 T�{w|7Bΐٱ��'���&��#�� �V��j
�H7?�Mo��^V��x�]b�q3(��H:����I��b�X�W}B�����h�X:�9P�ש�����cLApQy� ��I!kp��<�	�3����a�������6��#�'�O�N)Z(D/6>�D2�%P�3r��e�F���:缓F�s��N|�'��n�"]�]U�P�x1��i��^���F����6<��4+�#�í�Z?��v���J��V��ٌg���%���؃[����X�Ȏ]������-��I�����|���)c�_^C�=��~P߀��̺��c�K���eM	˗tp�d3{&��2$	&Ƴ
�ܿ:����ܬ�x�?�nn�
��V�z�X�@lӳ�G6��Yp�>���?o��Z���\��0-���"�l�|@�S�x��MږOq��i!T���o}h-\S.�4��b�[lT���	_\-,8��bܷ6��}ut����I�H�
9�iuk��R?��>ԊJ������C2��1�]JM^Y�sp�k�]�b�Śz>�b�s��������{ɒ����QP�󐌊�B��&Ix^S�0?� >
��@������-�h�FӺu��|�ǂ�5��^���m���.E+�G���#��I����ŀ�Nv�&�b�h�޳-B������e�Y��apvɾ����;�1R�g5B�I��U�Y���};um�}AP���ǚ~�c�Fr�+a��Ʌ*Щ������NNN��ds��]�A�ᨑ�פLo��)���/�yk��Om�`�o@�i�[��Fn���q��"�䨣��E~M�|��~qN=�=}W{����W�	���.y���U؀��P9+�W󉹗eA�Co0g�H�J�о]
�ܬ+�V\�)<������C�F�Z�hw�^>$Q8�4@�t ��A�ҞW���Z�~A����X{�|u���O�N	R��:���l�>='h@�7y�(!�'��&p���:��F	7��a��h̶2����C�ǟ�6�c����⌌R����+����r�A�U�u�-��Qp�!�5u�K[���TهK��}��1ߣ���&ֶ�`O�e������\�hty��Y���9&��w�S�*%���7�!|n�*m�&�k�_�<=�t�ث�Gմ�����t6]a�n�Y�S
A��^T�[�3���8Wn�,���ˌ��Y�\��;jW�X�?a9+�)��P��N	�)d,B6YG�]q�=ݼ@֚�(�"��Gs�q�oY��P�p�w@Ǆr��TP��p��FƘ�>>�~a�Nc\h�2
L?/X�������@���nr]��u���+�&�A�X����N��.M�K�����]0�߽���4O-E�៭-�z(�Ȓ�&�; / ����N�-&Uh���;j�������a�|j��ܬ����z�C	�s�jX�y��v��jQ${�W�2D�x���x�1-ڒ�<r�π�q�N��3�]�'���6B��?�/6d�x`����w���O�M��_������.V���Uf�$wL�$�ޮ��Rq-PP�������O&�28��6R��ڋ˅��v�M��ɂ��
wr��\�U6�C�-�Q�[(���4;hȩKI4A�A��GX7�>Ι�a�C�w {T-�f�� �f���P��{K4Ef���
�SC���cQ8�/�E�G�ο���!2?�c;���s:�L
���7��ʍ����m�"�?`̅��ZX��<�I#[�e.�������&�������Ex�o�����a�读!0	�H��W��}*5AI���>�TT��K:{����tU�ś�kZ��u��aϐ=�tU�7aB�do�Rˤ��	.�8����Pq��4<ПV�����~�����zal�F^�nvڣ�x ��q�l�,�Kq���$A����n�=�@�o�6!�/2\��H��H��&!꽓l�]0<�����)Ю���G9�\����J�ђÛ��%��k�V�p)j�`�ʉ��jB��i2�ѻإ�oE�M��*?E������f i�=��Fld q��H;��m�	�DPt�w�����nt�]����o�:`N������4���\ݩ�����9�(��u�������l��.|�`�E\b���Q��i�l�g��;��x�X�o�ߚ��^_	�h	�P�J�dN�-���!2�~�;>��+۾�i��E�z�R������:�q����<*:��0Q��+%aTfkB@U�'���j��w5V���c0�}��}<$��D2Vm4v��I��.%�kY���>���=U��U�;�\�����v�RI��Du�hM����rR�`����m�kZ,�����.�|7�볋Du˩n����}E�L�̠_8�����ۭ&���ұ���~����t���D؁b�#��0��M~��]�0��e�/�,��E���lIr}��s�+�C|��f��@�_��s�M��29��*M��Ո���&\D�[
��{>��Y�b;��]��68�RP��������ɖ�&��o��Q�}q�q�\�!a�yS��K}�K~�`ѵg�I�=��sN�|��.����Cڻ�x%�g,,*H�fw���ـ�h�"��[�pX��������jMV+`�e6���C�����l���e��f{ܯ���������,y�K�Zj�%F����>�7�.2(w�|Ԇht��T����bȫ7a��MC�J�q�`#�Q{0P�򽊿��|�Z�ݣ��]Q�v�O�]��8����
�ٿ��Y�i�����
 �Dƫ�����=��B�ݤ�Z��~���=8r�F���B��Ŏ��U���� ��6J���b��c!�*���{vDUha����L�u.�蔰px���ƉQ��@����eCˁ�:�~��@r������Ƴj
f���+νe���'[ �a���)��7ATt l��;�����"��P���*3 ���I����Ywc��-Fk��1yɿP=�z��������6vGolG~.�'�nn�x P�M%;H��aM2��y�Ӳ2�c�
��[<Z�ŝa�GRF��b�e��˛�VO�
�HL]~���N��ݞ�٩q؝.�y�{�K��W�:L������G�2�����I+�/v&��(���GހH-FDh0{3�Uu�_�xxY|��3�l��� �m�J��rZ��:M�����,�b��|@�����I��ũ�a,�ԣާ�[�)V'ʿr� &�-5��Ϭ� &>�F����8ȍ;.t[��Nj��o3 ��ʠ�.�
tMޖ�p��L`�g`���N�?�Qv��*�
WU��4D6�9Ɨ�Q�>�^���(�=�m	ǒ��(C}���x�ʜ�xU�h��F�g���h���`5��ބ�;]�o4y����?#ZU�������m��x�
pZ�l��:���,�T!��_Z��xW��1���������9��3,��ݾ��_������L�	�}�6V+e�1̊�L#�W�i+���d��߮��9OqH��'*}��&<����1{��VG}��"�ɨ|6t��A�䦘��pQTuG|"U�ɟ��!���,Wy�%���V^�W��o�4�/�]j	�ڜ�un%�.؉6ZB��zstئ�I[j/	���G��b$������B�1��!��U�c�Z�Ŋ�ǥ��:�ˌ�x!���Ұ��@�u��R-Pĉ_;�k*1���"���<Y��$��KНF�yMؑ��{��s�?(�y��>
�����c�%!�';�.�T��"g�5'F?�B��0��X�S�v�j�v�����#8�_:�.��� ����oc� >L������K<m9<�0�J�yi��;��S�*�K8�������i�$��;j2��&+����ЊD�޽"ΩV�9�J^��= p������x���O����\�uwe�ע��&�rA�֥z6>�_�������86w΄�[:�r�
�A9�=m�>�5w"R#����H��Es�$��?č؛N6�����7���~��� �F����"A0��,�e(xu���H뒋����60EKɏ3*5���Ô%&�����u�#������� l�0������}�Pȷ��Q�	�����œGkv��0Ǜ���`/x�,�zĈfu$�f(���s��2Q�d����J)��k���c��/qaErw�'�G�i�[���~�i���ʥ'��FB�ױ�������[�c	��e�J�3kg�j�@������>����M�h���/+�C�����Լk��7�.K��\9y�z&�����e�yw�5�(j:�;%I��%<�3�����́Ѕ���{K2���.�;���EvF��ȖMe�(�r�E���=��&�K�)���_��ٺ�d�C/��WJ$����X��/��r�C�r��R��y���"35��$��W<X��d���t���@XD�����"���I泞� %��lщ��K��)"�����$�C�
��A,:�Z��H06D�+�$�VLؠ����&g�$���Z�9��<Ln�F���m1�u�(�5�?�W���;*e�T���_^ܫR����HNm3���Al.%��ʀXTm��u�3{�ǩ��D�nԸ����	�1+y1�>:��g��V�k�sL��r�8|�&Y�����ٵ&��O}`��&7�K��"�d`�@�W���y8oF=�xmZ��Y�l�gf�b��<�$317�`֙J�mB�󰎮���]�;�HL-�<�o�%�Q�MqJ�H�ch�ˤ���((�\fu�[�-ɠ|6��)�t:���ޗ�P7���ܩ��p���8ZB�|�Z�0�!���11Ӗ'����_�L��4>�h)um	*'1��^�y}F�pø�����"c�P�� ^K7�"�m�y��lH%=0�� �ZI*�M����W/�id��L�?P9�)�1;nql��`�-�	�'���S�^1a�#q�ϥ�M�O1&y)T��3��guh W�s�:B:M=�uX]b's�"㦷�צU[ձ�f��uC�TI+I>���ll��uYSP�l�\��W�{��m�&]}�yc7խ;���} �|3�������y'�����a��_�~��U�����f9�=��s���z�Ԙ����3ٞ	��?�g�+o-���HP ����s�arf����g��:�M���]��+�{qt���������+�б�Ѐ�6�D���2*�:��5_�0[����"�HC�p�M7���j��G�v��ò�	7"� �HZ��J;��i��'�r���5B��ÁHF��$^�f�m�gy���kYf��7�b���M%�����r���婞GQ��NO��.8�@��AEi��*	i��V���Y��6���:9VpN�Ͱc����`��J��(�[�ı:�Fzn���������0�rI�
Ȼ�c�/b�[��	�cuYQy�P�D��e��*��Z�?k�=]20� 0�����%U��\��_�9xym��'��u97��BN*ѾGS�������L)٦s�gtk꼏e<;��^��l����nz?&H�DM�+۱(��6��R���/�SYMh���"!5�����gl����"����x�>���W53���uZ�(���Z�K�՚�J���uj���\ީ3��44� E�|�Q����Z]��݋��w�?���sf�1�K �u�:%V�>�Y�ҟs�;؅K�`�Q���J4?�<#8
�0F��4I�]۽JҲ^n�0>�t�ǰߛ��9���4$����fK��jZF����tp���s[�`�~���b�J�l�
	`��@Νh_;��8��-N{����iW^t���,
1��;������}(pp�-�Ӵ���w;��;S�~�|>`	� �����;,��2��ݔ��� ����;A��|���܁��Ň�4�:9�3����G���
kV��95h|�-3}����W������T��k���]�� ����Z?�]�A&�g������@@��Y�n7ڌ�o]�S��L�4��{0��ٮ�*��ND�I�m<DO+$I��4���X_�U�H�{�s9@�<��{VT����S���6����I��t�i��U^p��Џ<�2h_��C�Jlp�e�<B��ҦaB�������?��+�w�DțO�bb?�~�Pz���^���Γ�����'l���r��omG�5IuO)	��B�(e�}�.� ���s�����;<KBDr��caQ����]g��!̋� /eά%
ͱ����{-j�{�x��F�ǩt6�	=;J�hF|�jI�[E�1I$8]�H!�#�z9
5��NgE
�)%~��^c�s��<)��h,��]q�;uN\�XL7`G�k�=��i�M|D�O��_�Q�����5�; 𿭋><>��o�6)��Q�b�'��o�\u�~Q7���%����7H2$BS����G�G���G��h�W� �i�D�D�I�A.���C��'5Rr��5��e�~��/1>0�/���)MO�CR�����$,QAz$�5���l�a9ܱ�w����z .����_o�b� ���/��P�0l5�D�����sJ�8b ��e*F�V���@�gu9�if9�I.�����cƚ��*1<#�a~��E�����g\�(��WE����L�e�8�7j��ϩ���Ǯ����h��t(ǘ" ��Z���͂x(��[�B�)_ׅ��r�_e�R��M�/���E��z3�A6�H��YJn�ǵc�;K�D|����
U�hN���ߠHn)y�SxF1cB��(HQ��TR�����L��͗�x�.���,ð<(�i�0� 8U��Ԏ�â�ը�T���.�V��g�v(@CP���zٸ/���w�U9a�(Q�'欓��IQV[HȒP��Kg����tE]�����Ժi�vZ!AOyy
Ė�PA��JtSd�шQ��A��X��fz(}3z� <
x��ʘ�+�5�@�m����i���oF �KQ������������Ѻ����GY��Q�`4 ���4� 7;��0l�>B��x�~�d�c.�1�Dz��-�|�����%0̹�o]*���0b֔!��/�D��2@�s���d�罌�|`w�L�ؤt��&����^'�l��"��2\�C�G����`�j�H�C���#\�}�Ӵ�!��Q�^��� oje� �������9j(���2�[&��k��1H��k�Y����0�ւ*�餌l�	��aY�_��r$���/�c���Yz�����
��)2���"��&)�z��$���{��݆��?��[���<SH�O+Ϯ6���j$�[�N��q��B�'W��)������j�ќ7��3�6A�� �6uiI���.M�p��M���O��h�o%��\��,�@e���V����A�R�>!V�����RS�)6���.0g���L0S�&�r�}a�ca�1����������<��wR���nQKV���T�!{tuŗ��$��909���}r�j����A9�Y�'���?�=/�s�)g��	�k��Wh��߶��H�4&��n�|�Z��Y��G~l�y���e]$��7�Z�t�0ZJE���#��'�$��P�%����	T�����z�??�x��=�*�}�6>��*���¸��E%ެr��}D�`�@�ym^�ܩ��VWDے\�A�${�+���e��m���ݠQ���F��4#:�*��4r�[U��;�1��[7G��=\N��8�����>��|�q��屒`��⢱��6:�m��,ڳ��ʤ�Y� O
"U�;۴�y���tV/eu�A6�Kx��#̵�I�� 6ch�y��x2@��9Q�B��FovNаO�>\��kC���]���Zˌe��PL�I�qߎ�����Ą��R?�Tΰ����:�F�~�/'L�t��1M�%��҄��������1#��n8&(@�|aX�P��Z���.Wś8��ٽ �p�]���<{[�᭫�N�e��!��ۭj,|�]u*�ۋ���I��a��N�6�ǉ&|��va��\�>�+_Pd����^�Ȉ,F.Lk�������}���e0��p�xV�����=ki6��!P���<ɪJ̨)�8��;��԰#VO�Z�5}����`rl�k����9���d餟�װ�?eS��=Tg��$�
b�9W2��C$w�1�h���`��U$� �劥c����NAd�,���I0k1��m��QP�a��k�Pg��u��5�W��ۘ�m��o޶B!Z���lC$q�G�k0􆹎���?�S2�E��pՄ���!C��_^��\Ŋ?1�:�A���fu��R`=?�pZ4S�KBGr�3��ˌԴ���J��v��_���t��������>�&G���ly�ȭh�,�V��r�?;�NX����7T(�@�Gӻ�3�D����O�C�"��s�5��u?{m~�z�x�z�����P����������^S�n"T<0�n�3����Ji���o�5I���e���k|}� ��؀׌��0���Ykq����I	��Sx-�`����98@���u� ©{���K��9 ����o��6����ϡ��0��M2�otO������:�Ӂ]$�e�������@�F�j��As��@E�r�ؑE;<S�álP/!G(Veq�t�zq9]7n?�a	�BR�J�0��Q�E�-����ڱ�m*�@�)�����b*�:IV������I��!�o:D��=m�[��	����gM^E3W�;0_��E.^�cM}=�/
ړ¹���g�ϡ���g�s�5��_�}R
^hg��
���hE��)�	���������'_F�&^��#5��n9��l^��v�'��nk�sI����QC>�c�_��%�f~���'�mCs���L�KJ�(��$}Wr��!��wk> ��Rؗ�y=F'���[y�V��S5�.���﷑�͑�^#�����\[*�g���Ζ��A�-쩐�w�U��?���Τ�KˀA�L�=ǹ�3��ʜ�YV�v�\����]kO5�a���eE�N�։�)��Z��q�Cahi�t��
�JX�yI�<܅�������� 	�V���5Ҧ��=��S����3��	��t�bt��Y6�3P��������R��a*Oh2�7�E��Y�Å��D��Ï�Tݦ��lL�%�:w��L׳�3�j^�6,�c���к�*B�'xa�ƾ�:��3X�g54�Vr��*��o����d���y��RR�&�kά��&������6|}�C!��\��>�J�+0�/����y.�Q9����0="���D�U�KF�\,�rh�S20E�h���hh�D�7?b,���R'�Z�C�P�;� ��n�Z�k������N �1�.27�B���l]j��v�D���"X�g/_6/_g�0��V�]��é�]�NO�,�����a�gJ��j� ��PB�<�y������;rQ�8�"����!�˴������fLtN����/��T�:xW���UDu><v�#�T�ُ!!VK.D��D�6,߆@# ����IIG5� U���X<�h/W`i�d?��}�GlE*��Qb�7�O�����!r]���G�d��Gо���iCe%�rjS���mZ�_s��B2O�5O>��'R6N�YB��)��ؿn��ȷ>
Y�bT#��I��z����{\�Ǿd,���n�2hh���%� �zB�V�I�m7�
L��s�/n�
ļ�P;�@���ԧ!�_��O�5q��3Z�����!@2Vx �4'R���QEƴ�$��\��ʄ��5�v �u��m���.�Tz���ߖ��[��r�~c�`J`��a����[��ݲ����l5)���V8�dL���� 9`�&����%�R���2J�|v��S~ئZ�.���Y����{�7��y�dK߀\Y:2iU[��D'���lG4sS�|{��7{ѵ�� �g�D����)�1B.�X��[($�=�1)�[�D议-���<�f(�&j��7�p�|�4C��I�}�T3rQ���sV�/osW�]k�}!�C@Ab��o�Z���V:���:Ѡ�3s�I?z�-�V�\^�О0Q�F�6���nG��{��R��$���N���,��D�b�ٓ�m�qb���E��؛Q����͘����SQ�����{D�(�0��]�T'�2L(��-�)�imW�5G������Z8�[)���|0�_>�v��4�ӷ����9'!������)e��n�� }e/��n�t����?[�𾨷(+Kj: e��i�m�|�	h严C��'���sy�%�p��@����6��������>8��^����QI�E� 30唍�]ClP�h����[y01���AR0���
�q���5�*k� ��.ݞ��%��7����y�~�a�L����t-��\���!�ʇ��]��-�+���,�<�U�=�Y9nZ�3�����
�@�ά�#�k���:�F��D�F�-�� �Q����Ÿc�k��,8��o"<r��z���.�AA����L��r�(<��;R���p�():���I�Y3_��FIjŘ,���&��2	%b��2%y��y¬��������ќ�z<'��Gy�W���&��?%�oS�T���W�)���'fs�Z�U�o����io����� P�m�{�<�:��f�m��������~�N��At��5�8��r5'����~�&�9ˆ��0��y������^���6VT�A��:Q��3�m�y�ֲ(��C,�y��?xR�f��,왑�g�A�PV�*
3hx
�"���W8~��KV���94������<}~������:��*�V�>�L�;�\`*
c4Z�i���5����ΰl��Ho�]K��;���m*��7re�BljC2�ǭA�>*K&����Dsq�4C!�^=w}N`������V9'!>:6d\��ˮ��6p8|M��q5�o�z�_
�`2[�n%y��N�#��JaQ��,�Ȃ�҄�}�e3ӖU*�`���@ǈ���f���!9ay��}�m�D�Dl)0��JA�[Sޓē7+������j��+���R�p�ڶ����uj�ho+�S ɹ/q�������'��X��b�����J�G������)�J(q��r{b^����uޜD�g-y]`]���X,�� > �$��Py%���$�jt&���׷�gꟚ���S���[;:�������b��+����,�g�?�2��R��$^0=J��v�Л����P!�\���N�x�rT�F܂�;�Ȯ`�!5�=��p>���}v&�V["���T�5�;�;�ES��{�H`+se����^�c����vdܠA�-II�k;@��D���Ǝz��v�ǹ��\3PF�5���XLE b�͝���t��� f������+ .�i��G�y��0�Q���\p�@��ܰ�9��"�8d�����CVኢ�_]}q�)�.��x�$,�����ӓ&㈣L���IC`���:f��	"�?���+Z͖u���l���\�t|��)j���Q���䆮�-t�q#���[�}0���`=Y�ݫh���X	�ș�O����%+��N����h�{3 �'�f��d�D'��)�Q�Fӛ�j��~g�R�?+ �&K6��Z���*Lߐ����YcA̅7,�+���q'�م�,`�7���G8?�#^�>�~)4
Ak(A�K��7�z4,���o�>K����8Բwn�"k�0��� �(��y��'����v3a,�9<��EQ���.�"%��qd 	b���t*�x�	����ګϕ��j�y���.Y����/
0�'~nZ�*T���&,4ֺS^�l VA�@<m���z+� R��"%[��Yl�W�	(u�Ҕ����7A����AZA�Nñ��r|�s�ºd�������n��Pv[�B�,�~�.χ�',)�4�^n˚S�v�_��l{�p��p��,���5_�IOi+A� ��JF��ֈ���J��@���g
�P`�I�5��OoX���3��6"��&�N�PCeɈV_���Ԩ(<f�	�4�'[�/����D4P������/�ʧ��Vc��؎��ሔ���.������XAB�%q���	T-<�]�i~z�-��]5�[-��Jڈ�dRҫ�z�B3Ló�4�=�H��.2V˛����M'm�J	�MY{��_H��dkN��
Ȳ�'��y04<&Z06������'+�{i�	{L���֖��!�8�`$��������	���|;(�
���4}�I��i��wt,-h�n`��i�}���Q�Q�)�hif�T�0�] �8l�z�;P��#ۣK�N��`
�����۫^�IN%��`�SJ�鈟x/��w^��Q��Kc�bQЄy�32]��p��W.��̄%�ԥfH�yF�˲4�HP�!{��q������w�8YX�橿�oX3=u�sN,������'_��=^�:|y�W=8�,�Tt���H�J�}�7�
��\W1}{��S�c�Z�E��V\�Mͷe��;�*\խ����F2��}f3����RKR�H}�c�k����aL��v9�W7�L3I�jo�.��ʀ�90fUU�[й/��\`3�<����Qq�U�h��f ���-c�?�A�'.,�S��C�}:5/�mS$�\�ۘi�=f�����'�Q	��Z��%%��`_��\BQ e)A5 �ڟ۾͹�?�A��@{T����^s�]�Ar[��T�V��?��
��I���:���/tP������U c�����5"��=�,��=��d�ol^�Z��xr��L�r��n�m�aO
Rlښ� �a?���qD�'{)+�|��56��5��P�Y�G�ݟ��Q��<���s���{loH:��%y����_0��^d�̸sV݀�GY*)�4ՠ�e��p�-l+*���M	
�T�l��_��B����r`k���/����$��zY6��%�,5r�-?iv�de�9�5ϩ���Ɩ�w��[�$��i1�P::���AC�¢ ���A���\�_#�7��mȿ���6�"J#DG�N�$�����`)�>K�XY^���2��F�q��j�;NBR�oẉ�h�O��d Nh�摘�N���'M�0�	^�O$��{|�wt�8x᯶�������.޸�A�a�{�����ˈ��r74E��V��amd/(���h�_�%���ٌWWU��=�ʭ��|~* ˠ ����dg�ɳ2�aω���n4�MtV��v���p��kmn�j��R!3���Wx���x� ����
�S%8&㸶?���4�FGf������U��)Z�s��(@�-�M<U�/�F�@Fµ`Y���yQ�\�ޟ؃�Rб��������"/���eq�q �x�s�����x�^���3m���%�¦-_I��-��/��?,:�e�>�,,8MW1�u9�g ���� '-k��('��WySqI\G�~�9gG�w�9g!�L}���������	��}WS?j���\�)�٪ɢ��k��F�3l��U	'{�+�`�ͪ"�H޷~���K�8~R���ҡ�HK��X����R��R�:���?��@ϝ�(��f�R�!ŵp]����R>�>bm���ɓ�[��N11M��w[$�ƽe�lPП֞��&��l�@�_1�n��U��.Cy8\�y�i!���4ٗ��0Hh��H4⬐;���XP�{/y����H��s�����g��|��(�����/�x�m�^$E����l�¹*LBw���b�-a͡� ,#����=��b���|[n�B>���OP�tͷ)���8��BCc��RY�'�1&sہGs��e�kk�_�<i�� |�y���!��8�9��{�
zW� �z<� @����8A]��~���q_�.rt\Ȳ�\�,LN��ֽ$�X�ӔVᛃPѻ����	�1��P�tG:'v� �̯�z�쭯P��t@�d�_I��	4ŉla�7��v:��D�œ��%�g�fm[~��Lr*L���S�F~��B�_v��ߧ��߂��P59����@�S.����Ύd�����+,<&kьU}q�c�"]�T
 ��2w}j����hK�Y��7�q6X��\*jw_�bcP,��.(�����\QS���އ68 Q������!��5�{�|Ju%�c������7����
8�ϣ�}�J��3y�l��zt�9���jX�.ȷw�B3��9��ڵ�Mug�卄��3L�~���Ŋ6�ܺW���'t��F�:J?��}��=B�I��BW�R�#Z����r�r�O��G��,�}@0+�n��0	/���Q3�[��gLa#x���CM����l�齅�k��\N�����I���M��s��H�2Q�Y�����a<q��4�ۗ��O	��o���$����Y��H��R�r�
?O?��pn{��c�-�K�@�0��#��˻ �⇬�o�8��b���[��X�L�xW\739�k��� r*&5������,�j��P�	<�fQ:��t�z��t�U��hq�:���\\�Vdh}DD
�!�~�	2�Ψ;i���]���t���&֒��Ry��ju=}����0��|F�Ky*2���IzkҸ��f|J\)XU~��O�r��~�?��2�
���^��߇���O���tz�)�0���m_�#�ĒsD�1H��Z`�~5�%��ɕyM�go�v6y�����}y�-
��a2��F6�4�E�EDK����\��R�a#�I�Fl<����nP�E�.�圍8���Z��?R�y�9��}2֦�T�O�_%��Y  U�E�q��MiipMz�+���
�
L|��<�!��gU���n�v�Bvw�#.����b�hR����+��gf��>(Z���vČ�(�QP��g�I?�|i&F�\sb����A����Og>Y1�G�i~W/�/p�n������[�MQj]�[�1��::����'m�ȩh[n]��n.�����z�I�9:Ff�W󋦓ZW�M�$~h%�5?�IwO��[b�˅{����;�¾�0`fƱ��!��IX�^:��"{�NfO���!�I��������x�L����6vk����%��������$H���yE�};����D?��1��Ŏ�-�u3j���!!J:)C��-�	�S�J��3���bE8o������.�߱`��)!�#ocr���j<�)̴���v�C�l��1z$��pY��ɒO��\��J�^�v�ι{�g� [�Z?/ Hz,�F}�-���m���G���!�	7���>���ܸc�'���o=����������t^xKE�1�`�+�ߣ�ϫ;}us�	(�� ��T�c�'X\�l��п�!\UCq��;o��'B�s�܌ʞ.�#��	���p9���;Yе���?ѪP@�x?����2�@�8�vg��4-�h��a�Wn8�h�Lwec���sS��L�2�V�
Ix#w�	t�9PJs���0����hFڳ�L��[��c���SU��ē�fsGt ��R�f��k�Yn�z�U���t��]�#�T�]@I�
��V3J"Ni����1����S|H%uu�SE�J�����Ku�+��Sl�|�w�p��}��8T7�.��H�a,�ږ���
�gx[\J�����>5&��P�p �7���5D0K��ʜ-�'�f��R�Ԙj�^�$O�h��Ɖwi���-YO8b��g-h^�`����H�ȑ܁������Q�:._��RT�|^�>$�u@�R�+���H�H|y�$��lN���k�h��)WxWTx��g���Y}X�m�;�>r�"'�LO`6w���ۓI��cr�u������޹~ �JW�����+���Țu�8����/*����3b���;-�R����{�4��4�!"��k��mKũD0T�b�˅�@����\j��תe��̛m3i���(��5�69�8a�V�����\�9D��F�m��~�{�V��dv�kC�V�}���t��O�o1�~d��
�+(4`yc��|�gU�ʎ�-�t�}��Ds��r���һ�E:!e��^�V���P�opc�*�����N>[�\;
 ����(&9�	�_0E�v&��P}L�aہ�p�6����<D��a_�h���]15�OD)D�J�ڡ��Ӹ�z��I�E`�/^6��A�������W�Zn)�1�!��]���e�j�t"#(.qR��2��4Y�&�FItLq�ې���82�n߻K�oh5��p4h%�s 7K� h6鈃�VJ����J�3���	�z���$��1�\�h�Y�_��wGg$�#�vU�D�
X���k�+��%W�~�0&&�[͟.!EH`[�f�_ߒ�۹oKF��.}u�PbqH�$�Q��x�P��q��kq�"�
䃄ㅑ,�znY�f\��&1��v%�� �J"�q�^��L��6�Z)��������t���.���	��|� <Nz~�e冢��Ґԑ��|5f-
Ȫ�E���`?w�?@�zX� Xܰ��3��.:51n� 6	�Dn���#��Z�'k�3�Or~3�{�Gε�S|��n	�}#��@��y��v���/I�$>JD�A���_�G3�p���&��"��k<��� �L������M��ٌ-g�2_�9?�G��έ��cL��#0�!A�јiA���v{�&R!%xt0<d�1��r����0'Q֧W�,�v��2ߜl�ōc�B�u�=΂8;!?㤋�{��M������U��i�E���5�˪Œ�[��]��М���$���o�f	Y&`�����d��+=�Q״�W�*P]EF��̅d�V���lC�p� 'T2�X����d�L�A:�ћ$
�-N�/YQ&p]�4�J!\�����s�������o���K�h��ע:�61A��4���C�OƱIua����i��>�h�ntO��QnB���Y��a:�RkX�^����&i�k��nW�����C�{����w����VRxV�b�<֜g֪(,|��;BH�_�l��/BS�0X�%K��ЇRt�%#�^nH�דV/a��\d�Ȟ��)3s]<�͗#3�/#t��O������ʪ��Wh�z	n�o�L|���R3orxlq� ��+�1<�W��R�y�
��������XUO6Q$�����7O�ɉ�W�-*7{�1Ώ2���*����h���!q~�"�~ޓ���/�b��e�L��t_����hXL�#�d�2�Ba�9 $V3��0��1n#�	Q]�vEi��PP6�ݳM�юm! �˘�Z'����R�f�!/ծ�����z�4�;PH�#�wm�X�GoEG�ޥ���/�����QmY��C�*	��~Z�i��?����eH��3��Y�W4������S�e��I�B��1����@�$�Oѯi�x��P��C����&z�Oi� �_O����;��Z����-�W���"ԙQSO%��4��"����K;������wǴ��G�
]w�Tl8�= '->�=�+*Ҝx��f ����1����n���2ݞS @�aV�B��_�`�wm$h^hR#�長�"?N#���A����{,�ǽ�iq[Lާ��e�UO�Y�$��y��J��O|��tF�;�����������2,��p�.�3P-��b�?�dK��=f���zĄ�^�i8�DA�,�䙉��{���(�d����.�M��|]&��]<Mc�(���1Q�<�r���|~����4ol����M(��*���5�L�^�^C|3�57��5�@k�>b����O5���Yd�O�����^������Ͷ�0\��O�ir���sY\���d_�=���d,�����֩�Vԯ�c��z���Uq���B���	�c����V"(���Z��guF߶N�E^4�����r?
�=;�dq,MJ
���"�c��7�~kW�S��Z\����3! ��{g��f�ˀً��m��)sN��^�������a�h�ݮ�P F�x�1��\�\�fr�&�[
�L�A"����9�aGF�:	 t�"�Î�2��pF�ʶ"�āp��c��㹰U�)$]�����p�0F��c\K]�:Z�e�x��Df1�
f
�Gnظq(���0M���g�>
�?#��E�'��_0�k+�{�W�9Q'�&���01�U,+�m�#��-Ȍ�i§0/�T��eQ'�v}�@)�vlM��^���i΅q	����BnA�����/�W�^��T�%:��3�d�2=!�@^�i�XM��m)�s|�h+�q��*�rI6�b��Yzc�.*�}���=������#|�҃�f�`�07��%�x%���L��B�9��Y��:����[��6��o� �*s;p�(�m�#��k��	aj���!�Ǖ�DW�T]z&>��4�)�h/  �.���f~���֖��	��[l�<�+X9)�4o�&�7��aF38Z��S�{���w#�7>2%��K����K��5݅|�{�#j����4�7QE��,��A<:��U%�z�Xw[,���������d@�4��C|)߆%�ZgU&m)Rbn�y5ͳ�ɻ��d��H>>��V�p�j�j�o5�1������Y��*y�N�̒�~��>%#�?�&�w������J��D�ھ��"�X�T��^�7�p�@藜�v�TC�"~sH�-#6��y'���Bi�����	���t�қ���0)�����v^��� -A���&�r:���(��zD�<>CR�3���Z��g���ڼ��B�.9�[7+u�x~-���Q��`R�)��F����j����2�'������"]��Q%���5�B�t@�����w4�����0 e��S���>�ک�C�±(��H�k�<���_�q��L�6^��aC�ce�	}���aj(���CD-����	X�tx/�6��XE���ߪ��j�s�Py٬ȕ��p�0��̞ X]q�<4<�~ҫ}#��������p�8T��0���oq>�0l9�P��0���r�HK.-�k��@Ⱥ����y����'��kX�>�I�^�]e5���.�%�����`��h���w�����%����oU��!�����2cGz�E)�1D�!iPh���T! c�fT�4������{�¬o�P���x�@0�d-d�Zq�;,m��P���I�)	��,��h���)������^.��C�}N��c�U������D�W_���H�7jɪi��@U�"�0[p&zt3՞��Ƴ�-���� �N2��;��%��T�Ǟ���~O8q��.�+)5� �E������N��j��%�K��ьW:q�T���7,_KI_���;��6����%�0� ,?l����,S�;����D�f_;As����
A#�H/ܝ?�F��7�Ս���n?�3���?Wep)������R�A:�Md����=�1:�RQ��ɱ�y׌�������ȟh$�!�x��I��h5?��)��^�#4r��܆� ?\�׵��iiY��w�R��ĳQ���W�2A��q�d �[J��Ȗ�IdT���K��(�0?�C�2 �|5��T����#h%P�Hmh�=d�cc��Z�^����z���ro��k߆���W���]Fȃ�J{Oi��P�٠�@<Yk��������*�
�pv�^^,���=����2�!����γr�]�|M� 䈓�;�� ����!MZ��<z���r��T�\���j)�Մ���t�)%�*��n��*��\�.���#YI��.X}�{zn>VU4t�|�<���L�X[5.����u�����5��kV�c�\J×W[�
;�.�>�e�����:�����Q5N�AM�^���7���p42^9M��dy��Ꝭg�N��s��r��X��;&�k�LI󆷚�sk��h�$k��~�{B'[Q+^�����c��7Ӎ ������df�[��:��X�'�c��Y���c�ָ!����~�9��S�}&Ԅ��
��O'�0?]�
ߛ���ŚO�p�||B�r��emP�9���4��b��M������p/!�Ү�$0�c����h�uKh�KI� F�=��0��y��0������$�4����$}�L�{沮q9�@�|�T�W�ޙ�w#\+ ���L�n�����Ud_��չ~A�r�	��?}�|�O�<��������ݧ��$3#X)}&�uگn��懐���jACh�����?fP�?�[��&��A,����e���B윗��H8���q�к�F��A�|[>�����(�a-q�����Q���EYXC�˝���2�>XU�--�A)�w�;X�_�Yh���J]�-j�܂�ty�8
���tg��������: d���C�Q��W��a�L`µjq�1�ݬ��#�Q���[�-|�iQj!O��fD�_��d"a�I��N��P�(F�{m�w��?���
z�er�4�{�=���Ǻ��9��P��.p��߆�c��W� =�m�H�����$o� �韐�e�����D�Z��px��ɺ�Z�;�jSrt�:G����)���KFV����O���/�R���"" �b��z�dv,��R��|�Ek$�)K�? a�Q
��ޣc��!y������C�8z�F�A�� �Bx@��b�&OB6��m��������0�Tu�F�(��&�ug3��d���r�˦����Ot�)쉉���՟��;��@0��B��~Ӳb]ݺ��]6���/�ejߚ�Ǯ8�(B�E��@6�l.�X�t��6�Q>��Z�J��-�*���Z��j4��g_́�m���y��n�����B�E�+�i�l����	.�a���5�뜌c㓎ǟFz�±��A��9�R�3��
�K8��/�ȹ���f����q�����&��h��~9·�{���B��_�#MJl�v�
�#:Le���<*j��%���>+Kp�Yc�P�?��ۺ�N=�	/�C (h��ּл���ӳJɡ�
���p�/��U0G���}Tlq
���c�����+�ҫ��ۘ�5���@���h�#�;}�\�m�2
�Y��?�V/��8�AvP�˻� �X�EXrkI>##���NFQ,�P���dX����dN�T��NH�7�w*��QL�H��!u�t'��JX�b0vd��B�nY��0[q�q���[�t�Ea5R�4׋�p�"��_HJ�pJ3i�#u���T_���P��L�5pQV���Y.�7�.�`�1���o����(�����{���NMͿm��wg�쩹t��:�%�	�V�P��*9ٯ6�����'-Dn�����m����&�z�`mX�f�е�P����&0����F��XA>N}},.����f��	�?�����XO����o�k�j!�o/�{�a�w
����`��"�1�
SdY�ҟ�Fb%��J�_�}{]�[�>����ӳpoi��>�Y�꜄8d,�@�Ĭ~���xk���W����aO�v@���o����F� a�ė��(���w#�EB�<Ɇ�>�NIڏ��{��"��?�
&`�i-R�����8:��	�����j[Fډ�ݡ�L�x{� ����k[��F^�a�7��1Ă庇���Nv:f�q�ޣߛ]lC�f5%�k�P�K=�$+�.Fἂ3�p�T(d ���\��κ��%�V����#������&W�K��BsTyZ0�N�PE+�RW8��d�(P�uz�"�(���j�N��wE샡=�!qJ��sPy���Uh��'"��[a����|�����S�9�6D������iA��yx�
���T�ul �,����L�����ueȕ��bC<+}�$��8��Rf�b�Vx�
�2�*�2�vE/q�W��T��;��~�H�G�G^|	��J����|G�}W'�\?�:�6V�6�^���0����,�����\���Ig�-���e�U@~��>����bk�@5������Sa1"|K�Ns,�S��4�
̋n�"���=$>��GI�[�t��:
�x��Rz���#~�:����+Wmd���w�D5��y�J�y� �6	��߇7P�g�V�I6�<���Z"�0��c��0�����&+_uU1<_d���7�4���4�Hƾϗݖ�a}L�&�-`���Si��,�n��F>�⣹���8���ϯC�������80�ä3t�ezn)�xUD�Q�B�ElnhL�	(n4�cT��صL=�l+��� �PzL�a>����ᙨ����3��.�EB�y�,�ǭ����	��QG�vyOVC{`;8�	Ĳ������k�M* ����M�+�� _E{]@�������#P���T��*]�P�<}z��I6�Z�����Tѕ��ü	��׈��'y 3�P*�`3oPb@v5^��4fˍ)�����`���fG`%�/���Q�ݖz�W,��}O>�G���ɔ�^�"skZCԺ��9�tپJ������V����pc#�F�N@u�T�닶i
������'yE�i=�x�֯z�p�4Gfk)Mg���H�R\��#�6%����.�Y����jB��f��P�S�t�@'��8�f<�"�����hM�E�����K�s�2ܧۨS�1�ʐ�D�,?� x�o���Sαb^1*ȇ���\��4�`����Y�}��ڰ=C���qr�1�L��ޢQM)�0|!�+S�����:����hF�@(@���������E�#uާ��*U��/���^aq��ȡ����1�b��tD�zz�הC�
F�q�I�����nMv��d��\�E�^�<LB�x@`� �0��+N%�Ș�4���YLr�2�+Ct!�Cp7����Ͻ���Jt�I�� �J:w��n���Ac��j���Գ���݂�cu*�聩/�
�E���`�A��|���C��SFO��z||N���NA.y��8��W�W�s��`+�<l1,/h���X[�j�"�<��u	Z��׭x�T�o�C�s�o�����/������S�4���W
.���A�/�[�����۵G�c�/eL̀�.�.����<G��e>/�!�>A0w!�9�g�@s��dL@��`�({f�{rn�q�ֳg�v���y����b�?�QM�;wFj����#{2��%���W��T��KH&Ӻ ������A��*$�ɪ�c�o�P��xJ�Nb8۪P�"�8�Y-��S�ԲF��Q����h9x��AӐSp���y[g�VėȈ�R'GW�qAB�Ŵ�C�{��fFy�q�М��H��jD�I��0H@�Բ��超-��$Uu���(w��Kńi���N���jp< y֜i�ɶ6��qx� �h�y��_�o.�v���׭��T���	�Ҭ�9�MZ�Cb|L�����oڷ$B����ޢ}NI� 4@d_ogq�s��	�LV�S��r�z��Fd@�
	�
4G�xI���_1v$\a���s��5k7�D����r��r@?o!$7����Se�:�e���~�kBynR�� qi$�n��c���U8C	����!��4�+|L��[<���F�%�D�U]~��ю�������-��pb��$9#�Q��x	��LlY��)����H׾q���KK[��*,~�����c�t)��J�����n3ۤ�.��0�N��Yu�u�.~�����Y��f����>��1L������(y4���U��Ǆ�@v ���@���\��;�5��� �UBJC��p���,���.�ڦH4�����W.�m��@{a�8S�e���[���h��T+>�4&:�(���X�"e��tO����;j�˒/��G1I��;�n�cSFԧnqM%J�2��D�WR�$�8Va�6��;L�a�/�U�S��7��� +����8#s8TW^�g�m���zz;d�K����`X.s�8������݊((g
���y�}���^�R�&���,��Ǜ�8�?�_��Йr8��8ؑ�Q?�W)
̟��ۼC.��;c���z�?����9Q��^�tB���H�Y�R�=�!ѩo������a��A��9�f۸Nc�Y�>I�Q����a$�t��ii�Z�QnZA������H��d�}K��gZ^��Z���Tu��^o�7����I�k����}�,q�Z��<@ȭS�ln�O7��VC���AfT���񙎆_��ó�M�I��eU^fj������ 	��:F&>J�[HY��Q���;�R�M�����`0$,i��/P�p�%9���p�"bU�Qc�����u��� ��N	���;�/ͰR��u�F ]
�6� �覂^�I��4����=�ȊmJ��������NWkI�B ���~N5�M�l_w��{r����N?bu��RT�©�Dp.	�j���>������\����*����l�(4���N�kC;$h�����;-\�A��&h�F��ڠP�=�"���T��囏���'���aH�-rI�S�{��z����DK$F��2̮�Y6PMפL_�^r��-C8˗�#!{��.���9��^�k0����)�$��n��f�8��I��45>�5?��G761t�яg�v�l�p-K�Ĥ�/~SG�q�I�ެ
)�������~�4�D��>����z��JF���/욟���@�X+�ys^c����c�����\�0Q	�s��I��cܶ}PlC#��Go��~ui�w��M�8��n=�� �L �&Z�
�2c!1��&@2r����9�Y� �fn<2ō��]V��d�^����	p?a�+.��J��[��ƴ���. �b�����Qڱ\㵾�2>l�=)3�͸xQ�����d�&T���p9�:�;;�ʄ�:�=�
(�;� �K&+Q�;��͠� �<BH%A8�t��/����;z�*���Oί���}��
��`�p�� ��7�ߏ3/8;9D^��C�%�N��e��/�����AMDQb��rɀr���L��Z�닐��	��6��	��S����v�k�g�j�'�A�s�(�#��~�O�	F�Z�s	��)t�)����Hgǖ�����~�V�z=�
��Gzo��I[φ"O���_�����l�rT�@��spנ�LOog���!b��,�����J�x��(~ �;�|��n�ۮ;u��6�����e-��lŎ������iᤓ��H��γR�Iw��+UE�-<20*��� �M�v���l�>Ex>g^m����w�[�'���Z���K�S޼�d�E�6.�s���C��~C�)E�5I��W�؋��%/����Q��HÇ?���>�G;��%78G�F�ٽg,a��Lɯ:Q\19<�{�Pf#���9�����-v�T0/DG^,b#Ѕ��=fB]D��+Ą+W�� ~�n�2��M�p|N�j�V��y�&�4r8��e���Q�(�A1�7�<2��6�m;��+	Bc���o�����V����{\?/��d��W8�7�~����1pA�&�C�$��\����|����%!�����<�{��-�3���#U�jp+��3�c�;+X��>�~_g�K�lK����Ǯ^��Fc�{�֩��A&N��C�]#�:��P�dyz��gϹT��B�yE}Q�&�N��,yIl�0zP��J��K��P���u�^t���'r/�/�;��i~�\ �7#3o�\#(��i�=�2�H�Ŝ�>�I:�BP�6���f�{{��4�C�L^ }g�aո��K�a�hF����_v�|;]ƭI0�r��Q;$�ǝֹ��Q=@��=F�ӀK[p���
5{�c�G�렜d߱q	�D ����v�#��>����i�G���S��rz����q��&�<*젦���A�4� �+(dx����=���K�S,��g�6�y�[38'u��	�n�U)����Eh5j�� iF��h�Y+�7g	�ɹ6���=����-7�[gz=��0�b��j�Y�!Q.���A��*�)�(�y�9����j��<��!���7ѕ���T��e9U6
^lE�˒���pb��j�.�D���� $�`��?�p�u�^�}�g�@;X���}���q��];��X���D;ˑ�˔� �G����;]2Y/�-��^�5�5��ZuC�zd< �՚|�^�z(?��9i`���0�Sb͡�ԇ�,�V���/�-ޟ5�A��3�@W8,-��щ��;=����PBb�0ࠂcjЯ���BZ��h�&�alp��4�C��<�u�������<�7�)����P4���M�@ų�e�;vc���m\�e]g��ڐ���F��"�lҳ3w��-j���N3u;D(@Z��v_T�o}R��J�7�m(7V>/j|8/�(#

� */Uc~� 2w�g�� 7B�!1�O��5o������	W_%�>��,"_=�V��ھ�FTT�dV��Fv���Jo`��IK~����j2��	:*�c+n/����󃡖��ܤ�K�Ă�U�2��Y�)�>pҼDo�;�E$=���b'����=y�bvn��V��2��b^���`�[ل�g�ڻUg^8����E5�4
�}Ȟ���x��WN���F���ٔ��k��QmL���.��$��)�,y5��^���t�^̦���i��@�9���҉39�A��sXU�M�?"���&�ꓖˢeq���$�����j������j��Ti釻��5e���=���&LQ�'�|��aAqQ�������aZ5
Y �	�T{Jvר�eS۹	�U��
���j���ϛF���w������sr���'!�O���C�s~Mi-^�kG�O5s�`���h�Ju#G'����e�T��J�\��4�e$����A�d�̧cL�A_<3dt�"������yn�O�6��c-�g���O�	��ר^��ZMG����G5>�$�q0�J&M �HG�⠀�n�R�O�_�g����Kp�n��\ԡ��cX�ز���⧜Ђ�Yt�R 4!���N�����4�:��^���Yy?F���ZMT�;S��<�픸>U7�I�$�#?nW5��%�gK$R����:��?7�Y��PN|M��ON���K���b�Ј�C��Sq������2Y1o�� �ӤjD�;�J-���A�����m�GX�7�^
DK6������጗���縠�֧�'�P�_��],A�2���W/{+�S�hA�����j��?�Y�{�!�#�9�<�X�,�J1��G�v� ��_`����_���ks�QA,�H�ݟs��^�����0p�����N����&�Z���y�V�u/Y��<V�!ᰅ� ���n[n`**����KN� ]m-S@�AL7r�8(�=N�;Gu?�"Eq��U����Z���J�FdD���#?ۜT�,Ld�$�~.�ǁ�5�V�ذtenR���#��t9dO #��U�U�Q -tVl.��۠����p�	�n�8c���e�&-*i���U4^u��7L�US��>	�ځ�e���r�Jv��*+±ؠ����}��PA[i��3��꽥��� ��bA&m��T�
��)�����9g�YxiJ�jM{�z���0�L[b.�a��`���V�6B�o7� ،W�*����F%83�ث�Ō�k�Fu�)��*x�� ��&P��''�hш�M�[��a�Z��
���$O��ֱ��l|�j
�>ɆjD�]��#5�J�d6�����E6~8ȝP�qմR5W񏸘�]*�������z}�0*�l��/�I}M�5�l���4��d��0�}(��$�.�Y⩳������yQ��'�%2�n�~�E������ިy�P\P��"������%�H>�ové`���"�A �v|5�B����k��D S��f>(%��&����)��R~#`�d��d6Ш��ʨ{6��&�p&�^b��$�\P��$wP��M����fu+��#(�Q;՝[�إ�i��~���	���%�v��S�yR�#˱͍�ǎ�\��B��:����BNz��̅��E�����P�H�Pj��u-�,��,�3I�1g���ݢ2 N����uG�u,�S튤�n���d:���K��U]�$kb���,P�i��p�^u�
�Q`F_�2�4� �-nJ��)�(��� ��T�R��ZL�F��7����lr��^��,�&q�T����H+�% ���Qw�u?\��ɴ��Ob�dM�,�ʅB��]:����]�h2;���]�{�Ev9�H�A��B �AKH� M�PL@�o���9�K=�6-|��V�hN<��*�ls��?����=��2`�zh�8`o�#Ռ˧L c�B~h֌�d
 ��D�'��k�Kǘ29�����=�PE�_O)ː��OѩG5���J�©�cO}�)\F?c�C����8������:.�P�yG�8�i��c��)ӄ��Czl�oLVf(��s't�8��XR/�K]�7e���j���߱��=��w��ro'�ӧ�ۓ� *_�+>0�OT���vȢoK� �C�b�	m��Bbof�`Ì�i�A�K(h��H��V�ڭ��l�bd�A��
�IT�։+7�Oh�F�a�1J=k8���l���/j�1�����	ٮg����*"�D�=pJo��!l��+Ĳ���U���M�O������a^�>#���%�2X�?`[dV�9!V���?{,�AX"au��as�n�|gW�z�CR	ަ|0(�Q4�b"�l��A�CZ�ZY����uF�a��Y��Յ�XL+��?�(:B�_YU�吥��5�'�֢�s2E�E�c+��fI��!r�9O¥�[���7�ʔ�!�^��.l�xh�Q>�7�'2Ի���i�w�@����� �]&�q�&�~�֩>�?L�ԃzV����~"F0���:�)js��/L�}�_��x����v��ڢ��Y�I�zH�'����m^"qe�S�^�q�q���P`�����Bd�	){�JJ��ݘ����E�o��=�����|�i9�@��+���_�kB��~��{�!$�3F���H�ׁ�_�/��ޙ=�Q�/���d�܋^q�1POXZl�Iw��$�Q��-GB��}�)��$6��iAg@ߑ��fDC�����r�0�2�2���J#j���>����J�Mvh�J�9��D���&A�� @+�1���v����[��&�;���2���n�O�9�>�t�U)�Cb	�Xq�iIc��G���}S�{F����Ym%�o���v�-禛g�)���Wg��5J|�%��_+�ht+Hs+�@~ë(�ZJ��������F���(��}��PM�}:��K}�Vo?Dr�j��_l��L��e���LR��sQ��~��Bf�y��2�0�v��N\����ܔD��1k��f3�Ҳ�lr��ډ���ym�2�\�^(UF�K�:\�������Ȏ��!�f�5n)\�G�'���j$&�p����L ���8��f�F�5�A���([	�b��l~���S��rҲ�~�t
憈_��$cIgM�BBΥ��J�I���H,�&�w��>��G�|2>���h�+���	Ð�HkD�zk���T-,�l��C|�������P;&��;�T�|ZSy	&@Z�i�8^�~���:I�
�Q�ո_�?��RU|K!ע�9�>+��<�R�µ��_�7��q��Ջ�hV0|����"M��l�Cj�B���_l����x�ʶ>Iu�H���*������7t?�}���o��>=v��X�3+�W �	� ����6�~�+W��~��8J8����?���ޮׇ��,��ZR�n2D��+�c)�ؙ��_��-�[�I(�&|
��@���r�|V���޶*�*V��s���b�~��[%v `�c���L�vvh��}�g�,�JX���Dn~|��A���[�N�D:�#E����`Xj 0|澎F��s������M����*��iA �xe"��4�7I�(5v�\ny��S������Z�8J�-����^+�W��!���E��������T��b�����֖��B{����J#��EXz��nb�N�3�4��+��r�1�$K;�s���k�m��Ǟ���o�G�@���d߉dK�U��x<NZ�n��̐�[�����OV�w�ܲ�cA��/m����9_ѻ	������ֺ����T*ga�Ru��H�����������Om5	Xb��͂�۰�������.�Hp�⩵������9^�5��kN0����v��G�<�ݶI�||xJ 츮��a��%�I1~�I�ux�o�R�[�w&�>��.���IGA܉� P@��W�6�)fWHݽG�Lg��(���}|Ž�9B�<Ǭ�'���"�~Sevf3ط`�3Z��i��o��H#+�"��"��eaA�H+��o~py�^��zd��1�m����ߖ݉�6s��;j�̹��Bn#s��x��ֻHf)eޯxC1!��LN��|T�