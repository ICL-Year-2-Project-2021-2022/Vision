// Qsys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Qsys (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       //      alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,      //                                 .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                                 .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                                 .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                                 .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                                 .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                                 .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                                 .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                                 .vid_v
		input  wire        altpll_0_areset_conduit_export,            //          altpll_0_areset_conduit.export
		output wire        altpll_0_locked_conduit_export,            //          altpll_0_locked_conduit.export
		input  wire        clk_clk,                                   //                              clk.clk
		output wire        clk_sdram_clk,                             //                        clk_sdram.clk
		output wire        clk_vga_clk,                               //                          clk_vga.clk
		output wire        d8m_xclkin_clk,                            //                       d8m_xclkin.clk
		inout  wire        i2c_opencores_camera_export_scl_pad_io,    //      i2c_opencores_camera_export.scl_pad_io
		inout  wire        i2c_opencores_camera_export_sda_pad_io,    //                                 .sda_pad_io
		inout  wire        i2c_opencores_mipi_export_scl_pad_io,      //        i2c_opencores_mipi_export.scl_pad_io
		inout  wire        i2c_opencores_mipi_export_sda_pad_io,      //                                 .sda_pad_io
		input  wire [1:0]  key_external_connection_export,            //          key_external_connection.export
		output wire [9:0]  led_external_connection_export,            //          led_external_connection.export
		output wire        mipi_pwdn_n_external_connection_export,    //  mipi_pwdn_n_external_connection.export
		output wire        mipi_reset_n_external_connection_export,   // mipi_reset_n_external_connection.export
		input  wire        reset_reset_n,                             //                            reset.reset_n
		output wire [12:0] sdram_wire_addr,                           //                       sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                                 .ba
		output wire        sdram_wire_cas_n,                          //                                 .cas_n
		output wire        sdram_wire_cke,                            //                                 .cke
		output wire        sdram_wire_cs_n,                           //                                 .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                                 .dq
		output wire [1:0]  sdram_wire_dqm,                            //                                 .dqm
		output wire        sdram_wire_ras_n,                          //                                 .ras_n
		output wire        sdram_wire_we_n,                           //                                 .we_n
		input  wire [9:0]  sw_external_connection_export,             //           sw_external_connection.export
		input  wire        switch_export,                             //                           switch.export
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_sda,  //     terasic_auto_focus_0_conduit.vcm_i2c_sda
		input  wire        terasic_auto_focus_0_conduit_clk50,        //                                 .clk50
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_scl,  //                                 .vcm_i2c_scl
		input  wire [11:0] terasic_camera_0_conduit_end_D,            //     terasic_camera_0_conduit_end.D
		input  wire        terasic_camera_0_conduit_end_FVAL,         //                                 .FVAL
		input  wire        terasic_camera_0_conduit_end_LVAL,         //                                 .LVAL
		input  wire        terasic_camera_0_conduit_end_PIXCLK,       //                                 .PIXCLK
		input  wire        uart_0_rx_tx_rxd,                          //                     uart_0_rx_tx.rxd
		output wire        uart_0_rx_tx_txd                           //                                 .txd
	);

	wire         pixel_grabber_rgb_avalon_streaming_source_valid;                   // PIXEL_GRABBER_RGB:source_valid -> PIXEL_BUFFER_0:sink_valid
	wire  [23:0] pixel_grabber_rgb_avalon_streaming_source_data;                    // PIXEL_GRABBER_RGB:source_data -> PIXEL_BUFFER_0:sink_data
	wire         pixel_grabber_rgb_avalon_streaming_source_ready;                   // PIXEL_BUFFER_0:sink_ready -> PIXEL_GRABBER_RGB:source_ready
	wire         pixel_grabber_rgb_avalon_streaming_source_startofpacket;           // PIXEL_GRABBER_RGB:source_sop -> PIXEL_BUFFER_0:sink_sop
	wire         pixel_grabber_rgb_avalon_streaming_source_endofpacket;             // PIXEL_GRABBER_RGB:source_eop -> PIXEL_BUFFER_0:sink_eop
	wire         rgb_to_hsv_avalon_streaming_source_valid;                          // RGB_TO_HSV:source_valid -> PIXEL_GRABBER_HSV:sink_valid
	wire  [23:0] rgb_to_hsv_avalon_streaming_source_data;                           // RGB_TO_HSV:source_data -> PIXEL_GRABBER_HSV:sink_data
	wire         rgb_to_hsv_avalon_streaming_source_ready;                          // PIXEL_GRABBER_HSV:sink_ready -> RGB_TO_HSV:source_ready
	wire         rgb_to_hsv_avalon_streaming_source_startofpacket;                  // RGB_TO_HSV:source_sop -> PIXEL_GRABBER_HSV:sink_sop
	wire         rgb_to_hsv_avalon_streaming_source_endofpacket;                    // RGB_TO_HSV:source_eop -> PIXEL_GRABBER_HSV:sink_eop
	wire         pixel_grabber_hsv_avalon_streaming_source_valid;                   // PIXEL_GRABBER_HSV:source_valid -> COLOR_FILTER_0:sink_valid
	wire  [23:0] pixel_grabber_hsv_avalon_streaming_source_data;                    // PIXEL_GRABBER_HSV:source_data -> COLOR_FILTER_0:sink_data
	wire         pixel_grabber_hsv_avalon_streaming_source_ready;                   // COLOR_FILTER_0:sink_ready -> PIXEL_GRABBER_HSV:source_ready
	wire         pixel_grabber_hsv_avalon_streaming_source_startofpacket;           // PIXEL_GRABBER_HSV:source_sop -> COLOR_FILTER_0:sink_sop
	wire         pixel_grabber_hsv_avalon_streaming_source_endofpacket;             // PIXEL_GRABBER_HSV:source_eop -> COLOR_FILTER_0:sink_eop
	wire         com_counter_0_avalon_streaming_source_valid;                       // COM_COUNTER_0:source_valid -> EDGE_BINS_0:sink_valid
	wire  [23:0] com_counter_0_avalon_streaming_source_data;                        // COM_COUNTER_0:source_data -> EDGE_BINS_0:sink_data
	wire         com_counter_0_avalon_streaming_source_ready;                       // EDGE_BINS_0:sink_ready -> COM_COUNTER_0:source_ready
	wire         com_counter_0_avalon_streaming_source_startofpacket;               // COM_COUNTER_0:source_sop -> EDGE_BINS_0:sink_sop
	wire         com_counter_0_avalon_streaming_source_endofpacket;                 // COM_COUNTER_0:source_eop -> EDGE_BINS_0:sink_eop
	wire         edge_bins_0_avalon_streaming_source_valid;                         // EDGE_BINS_0:source_valid -> OBSTACLE_DIST_0:sink_valid
	wire  [23:0] edge_bins_0_avalon_streaming_source_data;                          // EDGE_BINS_0:source_data -> OBSTACLE_DIST_0:sink_data
	wire         edge_bins_0_avalon_streaming_source_ready;                         // OBSTACLE_DIST_0:sink_ready -> EDGE_BINS_0:source_ready
	wire         edge_bins_0_avalon_streaming_source_startofpacket;                 // EDGE_BINS_0:source_sop -> OBSTACLE_DIST_0:sink_sop
	wire         edge_bins_0_avalon_streaming_source_endofpacket;                   // EDGE_BINS_0:source_eop -> OBSTACLE_DIST_0:sink_eop
	wire         pixel_buffer_wb_0_avalon_streaming_source_valid;                   // PIXEL_BUFFER_WB_0:source_valid -> RGB_TO_HSV:sink_valid
	wire  [23:0] pixel_buffer_wb_0_avalon_streaming_source_data;                    // PIXEL_BUFFER_WB_0:source_data -> RGB_TO_HSV:sink_data
	wire         pixel_buffer_wb_0_avalon_streaming_source_ready;                   // RGB_TO_HSV:sink_ready -> PIXEL_BUFFER_WB_0:source_ready
	wire         pixel_buffer_wb_0_avalon_streaming_source_startofpacket;           // PIXEL_BUFFER_WB_0:source_sop -> RGB_TO_HSV:sink_sop
	wire         pixel_buffer_wb_0_avalon_streaming_source_endofpacket;             // PIXEL_BUFFER_WB_0:source_eop -> RGB_TO_HSV:sink_eop
	wire         terasic_camera_0_avalon_streaming_source_valid;                    // TERASIC_CAMERA_0:st_valid -> alt_vip_vfb_0:din_valid
	wire  [23:0] terasic_camera_0_avalon_streaming_source_data;                     // TERASIC_CAMERA_0:st_data -> alt_vip_vfb_0:din_data
	wire         terasic_camera_0_avalon_streaming_source_ready;                    // alt_vip_vfb_0:din_ready -> TERASIC_CAMERA_0:st_ready
	wire         terasic_camera_0_avalon_streaming_source_startofpacket;            // TERASIC_CAMERA_0:st_sop -> alt_vip_vfb_0:din_startofpacket
	wire         terasic_camera_0_avalon_streaming_source_endofpacket;              // TERASIC_CAMERA_0:st_eop -> alt_vip_vfb_0:din_endofpacket
	wire         color_filter_0_avalon_streaming_source_valid;                      // COLOR_FILTER_0:source_valid -> fir_0_0:din_valid
	wire  [23:0] color_filter_0_avalon_streaming_source_data;                       // COLOR_FILTER_0:source_data -> fir_0_0:din_data
	wire         color_filter_0_avalon_streaming_source_ready;                      // fir_0_0:din_ready -> COLOR_FILTER_0:source_ready
	wire         color_filter_0_avalon_streaming_source_startofpacket;              // COLOR_FILTER_0:source_sop -> fir_0_0:din_startofpacket
	wire         color_filter_0_avalon_streaming_source_endofpacket;                // COLOR_FILTER_0:source_eop -> fir_0_0:din_endofpacket
	wire         pixel_buffer_0_avalon_streaming_source_1_valid;                    // PIXEL_BUFFER_0:source_valid -> PIXEL_BUFFER_WB_0:sink_valid
	wire  [23:0] pixel_buffer_0_avalon_streaming_source_1_data;                     // PIXEL_BUFFER_0:source_data -> PIXEL_BUFFER_WB_0:sink_data
	wire         pixel_buffer_0_avalon_streaming_source_1_ready;                    // PIXEL_BUFFER_WB_0:sink_ready -> PIXEL_BUFFER_0:source_ready
	wire         pixel_buffer_0_avalon_streaming_source_1_startofpacket;            // PIXEL_BUFFER_0:source_sop -> PIXEL_BUFFER_WB_0:sink_sop
	wire         pixel_buffer_0_avalon_streaming_source_1_endofpacket;              // PIXEL_BUFFER_0:source_eop -> PIXEL_BUFFER_WB_0:sink_eop
	wire         fir_0_0_dout_valid;                                                // fir_0_0:dout_valid -> COM_COUNTER_0:sink_valid
	wire  [23:0] fir_0_0_dout_data;                                                 // fir_0_0:dout_data -> COM_COUNTER_0:sink_data
	wire         fir_0_0_dout_ready;                                                // COM_COUNTER_0:sink_ready -> fir_0_0:dout_ready
	wire         fir_0_0_dout_startofpacket;                                        // fir_0_0:dout_startofpacket -> COM_COUNTER_0:sink_sop
	wire         fir_0_0_dout_endofpacket;                                          // fir_0_0:dout_endofpacket -> COM_COUNTER_0:sink_eop
	wire         alt_vip_vfb_0_dout_valid;                                          // alt_vip_vfb_0:dout_valid -> TERASIC_AUTO_FOCUS_0:sink_valid
	wire  [23:0] alt_vip_vfb_0_dout_data;                                           // alt_vip_vfb_0:dout_data -> TERASIC_AUTO_FOCUS_0:sink_data
	wire         alt_vip_vfb_0_dout_ready;                                          // TERASIC_AUTO_FOCUS_0:sink_ready -> alt_vip_vfb_0:dout_ready
	wire         alt_vip_vfb_0_dout_startofpacket;                                  // alt_vip_vfb_0:dout_startofpacket -> TERASIC_AUTO_FOCUS_0:sink_sop
	wire         alt_vip_vfb_0_dout_endofpacket;                                    // alt_vip_vfb_0:dout_endofpacket -> TERASIC_AUTO_FOCUS_0:sink_eop
	wire         data_format_adapter_0_out_valid;                                   // data_format_adapter_0:out_valid -> alt_vip_itc_0:is_valid
	wire  [23:0] data_format_adapter_0_out_data;                                    // data_format_adapter_0:out_data -> alt_vip_itc_0:is_data
	wire         data_format_adapter_0_out_ready;                                   // alt_vip_itc_0:is_ready -> data_format_adapter_0:out_ready
	wire         data_format_adapter_0_out_startofpacket;                           // data_format_adapter_0:out_startofpacket -> alt_vip_itc_0:is_sop
	wire         data_format_adapter_0_out_endofpacket;                             // data_format_adapter_0:out_endofpacket -> alt_vip_itc_0:is_eop
	wire         altpll_2_c0_clk;                                                   // altpll_2:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, mm_interconnect_0:altpll_2_c0_clk, nios2_gen2:clk, onchip_memory2_0:clk, pio_0:clk, rst_controller_004:clk, rst_controller_005:clk, timer:clk, timer_0:clk, timer_1:clk]
	wire         altpll_1_c0_clk;                                                   // altpll_1:c0 -> [COLOR_FILTER_0:clk, COM_COUNTER_0:clk, EDGE_BINS_0:clk, OBSTACLE_DIST_0:clk, PIXEL_BUFFER_0:clk, PIXEL_BUFFER_WB_0:clk, PIXEL_GRABBER_HSV:clk, PIXEL_GRABBER_RGB:clk, RGB_TO_HSV:clk, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_002:in_clk_0_clk, dc_fifo_0:out_clk, dc_fifo_1:in_clk, fir_0_0:main_clock, mm_interconnect_0:altpll_1_c0_clk, rst_controller:clk]
	wire         altpll_0_c2_clk;                                                   // altpll_0:c2 -> [TERASIC_AUTO_FOCUS_0:clk, TERASIC_CAMERA_0:clk, alt_vip_itc_0:is_clk, alt_vip_vfb_0:clock, avalon_st_adapter_001:in_clk_0_clk, avalon_st_adapter_003:in_clk_0_clk, data_format_adapter_0:clk, dc_fifo_0:in_clk, dc_fifo_1:out_clk, mm_interconnect_0:altpll_0_c2_clk, mm_interconnect_1:altpll_0_c2_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_gen2_data_master_readdata;                                   // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                                // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                                // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [17:0] nios2_gen2_data_master_address;                                    // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                                 // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                       // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                              // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                                      // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                                  // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                            // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [17:0] nios2_gen2_instruction_master_address;                             // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                                // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_color_filter_0_avalon_mm_slave_chipselect;       // mm_interconnect_0:COLOR_FILTER_0_avalon_mm_slave_chipselect -> COLOR_FILTER_0:s_chipselect
	wire  [31:0] mm_interconnect_0_color_filter_0_avalon_mm_slave_readdata;         // COLOR_FILTER_0:s_readdata -> mm_interconnect_0:COLOR_FILTER_0_avalon_mm_slave_readdata
	wire   [3:0] mm_interconnect_0_color_filter_0_avalon_mm_slave_address;          // mm_interconnect_0:COLOR_FILTER_0_avalon_mm_slave_address -> COLOR_FILTER_0:s_address
	wire         mm_interconnect_0_color_filter_0_avalon_mm_slave_read;             // mm_interconnect_0:COLOR_FILTER_0_avalon_mm_slave_read -> COLOR_FILTER_0:s_read
	wire         mm_interconnect_0_color_filter_0_avalon_mm_slave_write;            // mm_interconnect_0:COLOR_FILTER_0_avalon_mm_slave_write -> COLOR_FILTER_0:s_write
	wire  [31:0] mm_interconnect_0_color_filter_0_avalon_mm_slave_writedata;        // mm_interconnect_0:COLOR_FILTER_0_avalon_mm_slave_writedata -> COLOR_FILTER_0:s_writedata
	wire         mm_interconnect_0_com_counter_0_avalon_mm_slave_chipselect;        // mm_interconnect_0:COM_COUNTER_0_avalon_mm_slave_chipselect -> COM_COUNTER_0:s_chipselect
	wire  [31:0] mm_interconnect_0_com_counter_0_avalon_mm_slave_readdata;          // COM_COUNTER_0:s_readdata -> mm_interconnect_0:COM_COUNTER_0_avalon_mm_slave_readdata
	wire   [3:0] mm_interconnect_0_com_counter_0_avalon_mm_slave_address;           // mm_interconnect_0:COM_COUNTER_0_avalon_mm_slave_address -> COM_COUNTER_0:s_address
	wire         mm_interconnect_0_com_counter_0_avalon_mm_slave_read;              // mm_interconnect_0:COM_COUNTER_0_avalon_mm_slave_read -> COM_COUNTER_0:s_read
	wire         mm_interconnect_0_com_counter_0_avalon_mm_slave_write;             // mm_interconnect_0:COM_COUNTER_0_avalon_mm_slave_write -> COM_COUNTER_0:s_write
	wire  [31:0] mm_interconnect_0_com_counter_0_avalon_mm_slave_writedata;         // mm_interconnect_0:COM_COUNTER_0_avalon_mm_slave_writedata -> COM_COUNTER_0:s_writedata
	wire         mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_chipselect;           // mm_interconnect_0:RGB_TO_HSV_avalon_mm_slave_chipselect -> RGB_TO_HSV:s_chipselect
	wire  [31:0] mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_readdata;             // RGB_TO_HSV:s_readdata -> mm_interconnect_0:RGB_TO_HSV_avalon_mm_slave_readdata
	wire   [3:0] mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_address;              // mm_interconnect_0:RGB_TO_HSV_avalon_mm_slave_address -> RGB_TO_HSV:s_address
	wire         mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_read;                 // mm_interconnect_0:RGB_TO_HSV_avalon_mm_slave_read -> RGB_TO_HSV:s_read
	wire         mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_write;                // mm_interconnect_0:RGB_TO_HSV_avalon_mm_slave_write -> RGB_TO_HSV:s_write
	wire  [31:0] mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_writedata;            // mm_interconnect_0:RGB_TO_HSV_avalon_mm_slave_writedata -> RGB_TO_HSV:s_writedata
	wire         mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_chipselect;    // mm_interconnect_0:PIXEL_GRABBER_RGB_avalon_mm_slave_chipselect -> PIXEL_GRABBER_RGB:s_chipselect
	wire  [31:0] mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_readdata;      // PIXEL_GRABBER_RGB:s_readdata -> mm_interconnect_0:PIXEL_GRABBER_RGB_avalon_mm_slave_readdata
	wire   [3:0] mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_address;       // mm_interconnect_0:PIXEL_GRABBER_RGB_avalon_mm_slave_address -> PIXEL_GRABBER_RGB:s_address
	wire         mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_read;          // mm_interconnect_0:PIXEL_GRABBER_RGB_avalon_mm_slave_read -> PIXEL_GRABBER_RGB:s_read
	wire         mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_write;         // mm_interconnect_0:PIXEL_GRABBER_RGB_avalon_mm_slave_write -> PIXEL_GRABBER_RGB:s_write
	wire  [31:0] mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_writedata;     // mm_interconnect_0:PIXEL_GRABBER_RGB_avalon_mm_slave_writedata -> PIXEL_GRABBER_RGB:s_writedata
	wire         mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_chipselect;    // mm_interconnect_0:PIXEL_GRABBER_HSV_avalon_mm_slave_chipselect -> PIXEL_GRABBER_HSV:s_chipselect
	wire  [31:0] mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_readdata;      // PIXEL_GRABBER_HSV:s_readdata -> mm_interconnect_0:PIXEL_GRABBER_HSV_avalon_mm_slave_readdata
	wire   [3:0] mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_address;       // mm_interconnect_0:PIXEL_GRABBER_HSV_avalon_mm_slave_address -> PIXEL_GRABBER_HSV:s_address
	wire         mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_read;          // mm_interconnect_0:PIXEL_GRABBER_HSV_avalon_mm_slave_read -> PIXEL_GRABBER_HSV:s_read
	wire         mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_write;         // mm_interconnect_0:PIXEL_GRABBER_HSV_avalon_mm_slave_write -> PIXEL_GRABBER_HSV:s_write
	wire  [31:0] mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_writedata;     // mm_interconnect_0:PIXEL_GRABBER_HSV_avalon_mm_slave_writedata -> PIXEL_GRABBER_HSV:s_writedata
	wire         mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_chipselect;       // mm_interconnect_0:PIXEL_BUFFER_0_avalon_mm_slave_chipselect -> PIXEL_BUFFER_0:s_chipselect
	wire  [31:0] mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_readdata;         // PIXEL_BUFFER_0:s_readdata -> mm_interconnect_0:PIXEL_BUFFER_0_avalon_mm_slave_readdata
	wire  [13:0] mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_address;          // mm_interconnect_0:PIXEL_BUFFER_0_avalon_mm_slave_address -> PIXEL_BUFFER_0:s_address
	wire         mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_read;             // mm_interconnect_0:PIXEL_BUFFER_0_avalon_mm_slave_read -> PIXEL_BUFFER_0:s_read
	wire         mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_write;            // mm_interconnect_0:PIXEL_BUFFER_0_avalon_mm_slave_write -> PIXEL_BUFFER_0:s_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_writedata;        // mm_interconnect_0:PIXEL_BUFFER_0_avalon_mm_slave_writedata -> PIXEL_BUFFER_0:s_writedata
	wire         mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_chipselect;      // mm_interconnect_0:OBSTACLE_DIST_0_avalon_mm_slave_chipselect -> OBSTACLE_DIST_0:s_chipselect
	wire  [31:0] mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_readdata;        // OBSTACLE_DIST_0:s_readdata -> mm_interconnect_0:OBSTACLE_DIST_0_avalon_mm_slave_readdata
	wire   [3:0] mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_address;         // mm_interconnect_0:OBSTACLE_DIST_0_avalon_mm_slave_address -> OBSTACLE_DIST_0:s_address
	wire         mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_read;            // mm_interconnect_0:OBSTACLE_DIST_0_avalon_mm_slave_read -> OBSTACLE_DIST_0:s_read
	wire         mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_write;           // mm_interconnect_0:OBSTACLE_DIST_0_avalon_mm_slave_write -> OBSTACLE_DIST_0:s_write
	wire  [31:0] mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_writedata;       // mm_interconnect_0:OBSTACLE_DIST_0_avalon_mm_slave_writedata -> OBSTACLE_DIST_0:s_writedata
	wire         mm_interconnect_0_edge_bins_0_avalon_mm_slave_chipselect;          // mm_interconnect_0:EDGE_BINS_0_avalon_mm_slave_chipselect -> EDGE_BINS_0:s_chipselect
	wire  [31:0] mm_interconnect_0_edge_bins_0_avalon_mm_slave_readdata;            // EDGE_BINS_0:s_readdata -> mm_interconnect_0:EDGE_BINS_0_avalon_mm_slave_readdata
	wire   [4:0] mm_interconnect_0_edge_bins_0_avalon_mm_slave_address;             // mm_interconnect_0:EDGE_BINS_0_avalon_mm_slave_address -> EDGE_BINS_0:s_address
	wire         mm_interconnect_0_edge_bins_0_avalon_mm_slave_read;                // mm_interconnect_0:EDGE_BINS_0_avalon_mm_slave_read -> EDGE_BINS_0:s_read
	wire         mm_interconnect_0_edge_bins_0_avalon_mm_slave_write;               // mm_interconnect_0:EDGE_BINS_0_avalon_mm_slave_write -> EDGE_BINS_0:s_write
	wire  [31:0] mm_interconnect_0_edge_bins_0_avalon_mm_slave_writedata;           // mm_interconnect_0:EDGE_BINS_0_avalon_mm_slave_writedata -> EDGE_BINS_0:s_writedata
	wire         mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_chipselect;    // mm_interconnect_0:PIXEL_BUFFER_WB_0_avalon_mm_slave_chipselect -> PIXEL_BUFFER_WB_0:s_chipselect
	wire  [31:0] mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_readdata;      // PIXEL_BUFFER_WB_0:s_readdata -> mm_interconnect_0:PIXEL_BUFFER_WB_0_avalon_mm_slave_readdata
	wire   [8:0] mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_address;       // mm_interconnect_0:PIXEL_BUFFER_WB_0_avalon_mm_slave_address -> PIXEL_BUFFER_WB_0:s_address
	wire         mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_read;          // mm_interconnect_0:PIXEL_BUFFER_WB_0_avalon_mm_slave_read -> PIXEL_BUFFER_WB_0:s_read
	wire         mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_write;         // mm_interconnect_0:PIXEL_BUFFER_WB_0_avalon_mm_slave_write -> PIXEL_BUFFER_WB_0:s_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_writedata;     // mm_interconnect_0:PIXEL_BUFFER_WB_0_avalon_mm_slave_writedata -> PIXEL_BUFFER_WB_0:s_writedata
	wire         mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect;    // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_chipselect -> i2c_opencores_mipi:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata;      // i2c_opencores_mipi:wb_dat_o -> mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest;   // i2c_opencores_mipi:wb_ack_o -> mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address;       // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_address -> i2c_opencores_mipi:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write;         // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_write -> i2c_opencores_mipi:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata;     // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_writedata -> i2c_opencores_mipi:wb_dat_i
	wire         mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect;  // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_chipselect -> i2c_opencores_camera:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata;    // i2c_opencores_camera:wb_dat_o -> mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest; // i2c_opencores_camera:wb_ack_o -> mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address;     // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_address -> i2c_opencores_camera:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write;       // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_write -> i2c_opencores_camera:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata;   // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_writedata -> i2c_opencores_camera:wb_dat_i
	wire  [31:0] mm_interconnect_0_fir_0_0_control_readdata;                        // fir_0_0:control_readdata -> mm_interconnect_0:fir_0_0_control_readdata
	wire         mm_interconnect_0_fir_0_0_control_waitrequest;                     // fir_0_0:control_waitrequest -> mm_interconnect_0:fir_0_0_control_waitrequest
	wire   [8:0] mm_interconnect_0_fir_0_0_control_address;                         // mm_interconnect_0:fir_0_0_control_address -> fir_0_0:control_address
	wire         mm_interconnect_0_fir_0_0_control_read;                            // mm_interconnect_0:fir_0_0_control_read -> fir_0_0:control_read
	wire   [3:0] mm_interconnect_0_fir_0_0_control_byteenable;                      // mm_interconnect_0:fir_0_0_control_byteenable -> fir_0_0:control_byteenable
	wire         mm_interconnect_0_fir_0_0_control_readdatavalid;                   // fir_0_0:control_readdatavalid -> mm_interconnect_0:fir_0_0_control_readdatavalid
	wire         mm_interconnect_0_fir_0_0_control_write;                           // mm_interconnect_0:fir_0_0_control_write -> fir_0_0:control_write
	wire  [31:0] mm_interconnect_0_fir_0_0_control_writedata;                       // mm_interconnect_0:fir_0_0_control_writedata -> fir_0_0:control_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;               // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;             // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;          // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;          // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;              // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                 // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;                // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;            // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire         mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect;         // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect -> TERASIC_AUTO_FOCUS_0:s_chipselect
	wire  [31:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata;           // TERASIC_AUTO_FOCUS_0:s_readdata -> mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata
	wire   [2:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address;            // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_address -> TERASIC_AUTO_FOCUS_0:s_address
	wire         mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read;               // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_read -> TERASIC_AUTO_FOCUS_0:s_read
	wire         mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write;              // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_write -> TERASIC_AUTO_FOCUS_0:s_write
	wire  [31:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata;          // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata -> TERASIC_AUTO_FOCUS_0:s_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                     // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                      // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                         // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                        // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                    // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_altpll_1_pll_slave_readdata;                     // altpll_1:readdata -> mm_interconnect_0:altpll_1_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_1_pll_slave_address;                      // mm_interconnect_0:altpll_1_pll_slave_address -> altpll_1:address
	wire         mm_interconnect_0_altpll_1_pll_slave_read;                         // mm_interconnect_0:altpll_1_pll_slave_read -> altpll_1:read
	wire         mm_interconnect_0_altpll_1_pll_slave_write;                        // mm_interconnect_0:altpll_1_pll_slave_write -> altpll_1:write
	wire  [31:0] mm_interconnect_0_altpll_1_pll_slave_writedata;                    // mm_interconnect_0:altpll_1_pll_slave_writedata -> altpll_1:writedata
	wire  [31:0] mm_interconnect_0_altpll_2_pll_slave_readdata;                     // altpll_2:readdata -> mm_interconnect_0:altpll_2_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_2_pll_slave_address;                      // mm_interconnect_0:altpll_2_pll_slave_address -> altpll_2:address
	wire         mm_interconnect_0_altpll_2_pll_slave_read;                         // mm_interconnect_0:altpll_2_pll_slave_read -> altpll_2:read
	wire         mm_interconnect_0_altpll_2_pll_slave_write;                        // mm_interconnect_0:altpll_2_pll_slave_write -> altpll_2:write
	wire  [31:0] mm_interconnect_0_altpll_2_pll_slave_writedata;                    // mm_interconnect_0:altpll_2_pll_slave_writedata -> altpll_2:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                  // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                    // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;                     // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                  // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                       // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                   // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                       // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                             // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                               // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                  // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                              // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                               // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                 // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                  // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                                    // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                  // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                                   // mm_interconnect_0:sw_s1_address -> sw:address
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                 // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                  // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_mipi_reset_n_s1_chipselect;                      // mm_interconnect_0:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire  [31:0] mm_interconnect_0_mipi_reset_n_s1_readdata;                        // mipi_reset_n:readdata -> mm_interconnect_0:mipi_reset_n_s1_readdata
	wire   [1:0] mm_interconnect_0_mipi_reset_n_s1_address;                         // mm_interconnect_0:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire         mm_interconnect_0_mipi_reset_n_s1_write;                           // mm_interconnect_0:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire  [31:0] mm_interconnect_0_mipi_reset_n_s1_writedata;                       // mm_interconnect_0:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire         mm_interconnect_0_mipi_pwdn_n_s1_chipselect;                       // mm_interconnect_0:mipi_pwdn_n_s1_chipselect -> mipi_pwdn_n:chipselect
	wire  [31:0] mm_interconnect_0_mipi_pwdn_n_s1_readdata;                         // mipi_pwdn_n:readdata -> mm_interconnect_0:mipi_pwdn_n_s1_readdata
	wire   [1:0] mm_interconnect_0_mipi_pwdn_n_s1_address;                          // mm_interconnect_0:mipi_pwdn_n_s1_address -> mipi_pwdn_n:address
	wire         mm_interconnect_0_mipi_pwdn_n_s1_write;                            // mm_interconnect_0:mipi_pwdn_n_s1_write -> mipi_pwdn_n:write_n
	wire  [31:0] mm_interconnect_0_mipi_pwdn_n_s1_writedata;                        // mm_interconnect_0:mipi_pwdn_n_s1_writedata -> mipi_pwdn_n:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                            // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                              // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                               // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                  // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                         // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                 // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                             // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                           // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                             // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                              // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                            // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect;                             // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                               // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                                // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                                  // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                              // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                           // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                             // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                              // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                            // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         alt_vip_vfb_0_read_master_waitrequest;                             // mm_interconnect_1:alt_vip_vfb_0_read_master_waitrequest -> alt_vip_vfb_0:read_master_av_waitrequest
	wire  [31:0] alt_vip_vfb_0_read_master_readdata;                                // mm_interconnect_1:alt_vip_vfb_0_read_master_readdata -> alt_vip_vfb_0:read_master_av_readdata
	wire  [31:0] alt_vip_vfb_0_read_master_address;                                 // alt_vip_vfb_0:read_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_read_master_address
	wire         alt_vip_vfb_0_read_master_read;                                    // alt_vip_vfb_0:read_master_av_read -> mm_interconnect_1:alt_vip_vfb_0_read_master_read
	wire         alt_vip_vfb_0_read_master_readdatavalid;                           // mm_interconnect_1:alt_vip_vfb_0_read_master_readdatavalid -> alt_vip_vfb_0:read_master_av_readdatavalid
	wire   [2:0] alt_vip_vfb_0_read_master_burstcount;                              // alt_vip_vfb_0:read_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_read_master_burstcount
	wire         alt_vip_vfb_0_write_master_waitrequest;                            // mm_interconnect_1:alt_vip_vfb_0_write_master_waitrequest -> alt_vip_vfb_0:write_master_av_waitrequest
	wire  [31:0] alt_vip_vfb_0_write_master_address;                                // alt_vip_vfb_0:write_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_write_master_address
	wire         alt_vip_vfb_0_write_master_write;                                  // alt_vip_vfb_0:write_master_av_write -> mm_interconnect_1:alt_vip_vfb_0_write_master_write
	wire  [31:0] alt_vip_vfb_0_write_master_writedata;                              // alt_vip_vfb_0:write_master_av_writedata -> mm_interconnect_1:alt_vip_vfb_0_write_master_writedata
	wire   [2:0] alt_vip_vfb_0_write_master_burstcount;                             // alt_vip_vfb_0:write_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_write_master_burstcount
	wire         mm_interconnect_1_sdram_s1_chipselect;                             // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_1_sdram_s1_readdata;                               // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire         mm_interconnect_1_sdram_s1_waitrequest;                            // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_1_sdram_s1_address;                                // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_1_sdram_s1_read;                                   // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_1_sdram_s1_byteenable;                             // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_1_sdram_s1_readdatavalid;                          // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire         mm_interconnect_1_sdram_s1_write;                                  // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_1_sdram_s1_writedata;                              // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire         irq_mapper_receiver3_irq;                                          // timer:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver5_irq;                                          // timer_0:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                          // pio_0:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                          // timer_1:irq -> irq_mapper:receiver7_irq
	wire  [31:0] nios2_gen2_irq_irq;                                                // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         irq_mapper_receiver0_irq;                                          // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                     // i2c_opencores_mipi:wb_inta_o -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                          // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                 // i2c_opencores_camera:wb_inta_o -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                          // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                 // jtag_uart:av_irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver4_irq;                                          // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                 // uart_0:irq -> irq_synchronizer_003:receiver_irq
	wire         obstacle_dist_0_avalon_streaming_source_valid;                     // OBSTACLE_DIST_0:source_valid -> avalon_st_adapter:in_0_valid
	wire  [23:0] obstacle_dist_0_avalon_streaming_source_data;                      // OBSTACLE_DIST_0:source_data -> avalon_st_adapter:in_0_data
	wire         obstacle_dist_0_avalon_streaming_source_ready;                     // avalon_st_adapter:in_0_ready -> OBSTACLE_DIST_0:source_ready
	wire         obstacle_dist_0_avalon_streaming_source_startofpacket;             // OBSTACLE_DIST_0:source_sop -> avalon_st_adapter:in_0_startofpacket
	wire         obstacle_dist_0_avalon_streaming_source_endofpacket;               // OBSTACLE_DIST_0:source_eop -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                     // avalon_st_adapter:out_0_valid -> dc_fifo_1:in_valid
	wire  [23:0] avalon_st_adapter_out_0_data;                                      // avalon_st_adapter:out_0_data -> dc_fifo_1:in_data
	wire         avalon_st_adapter_out_0_ready;                                     // dc_fifo_1:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                             // avalon_st_adapter:out_0_startofpacket -> dc_fifo_1:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                               // avalon_st_adapter:out_0_endofpacket -> dc_fifo_1:in_endofpacket
	wire   [1:0] avalon_st_adapter_out_0_empty;                                     // avalon_st_adapter:out_0_empty -> dc_fifo_1:in_empty
	wire         terasic_auto_focus_0_dout_valid;                                   // TERASIC_AUTO_FOCUS_0:source_valid -> avalon_st_adapter_001:in_0_valid
	wire  [23:0] terasic_auto_focus_0_dout_data;                                    // TERASIC_AUTO_FOCUS_0:source_data -> avalon_st_adapter_001:in_0_data
	wire         terasic_auto_focus_0_dout_ready;                                   // avalon_st_adapter_001:in_0_ready -> TERASIC_AUTO_FOCUS_0:source_ready
	wire         terasic_auto_focus_0_dout_startofpacket;                           // TERASIC_AUTO_FOCUS_0:source_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire         terasic_auto_focus_0_dout_endofpacket;                             // TERASIC_AUTO_FOCUS_0:source_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;                                 // avalon_st_adapter_001:out_0_valid -> dc_fifo_0:in_valid
	wire  [23:0] avalon_st_adapter_001_out_0_data;                                  // avalon_st_adapter_001:out_0_data -> dc_fifo_0:in_data
	wire         avalon_st_adapter_001_out_0_ready;                                 // dc_fifo_0:in_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;                         // avalon_st_adapter_001:out_0_startofpacket -> dc_fifo_0:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                           // avalon_st_adapter_001:out_0_endofpacket -> dc_fifo_0:in_endofpacket
	wire   [1:0] avalon_st_adapter_001_out_0_empty;                                 // avalon_st_adapter_001:out_0_empty -> dc_fifo_0:in_empty
	wire         dc_fifo_0_out_valid;                                               // dc_fifo_0:out_valid -> avalon_st_adapter_002:in_0_valid
	wire  [23:0] dc_fifo_0_out_data;                                                // dc_fifo_0:out_data -> avalon_st_adapter_002:in_0_data
	wire         dc_fifo_0_out_ready;                                               // avalon_st_adapter_002:in_0_ready -> dc_fifo_0:out_ready
	wire         dc_fifo_0_out_startofpacket;                                       // dc_fifo_0:out_startofpacket -> avalon_st_adapter_002:in_0_startofpacket
	wire         dc_fifo_0_out_endofpacket;                                         // dc_fifo_0:out_endofpacket -> avalon_st_adapter_002:in_0_endofpacket
	wire   [1:0] dc_fifo_0_out_empty;                                               // dc_fifo_0:out_empty -> avalon_st_adapter_002:in_0_empty
	wire         avalon_st_adapter_002_out_0_valid;                                 // avalon_st_adapter_002:out_0_valid -> PIXEL_GRABBER_RGB:sink_valid
	wire  [23:0] avalon_st_adapter_002_out_0_data;                                  // avalon_st_adapter_002:out_0_data -> PIXEL_GRABBER_RGB:sink_data
	wire         avalon_st_adapter_002_out_0_ready;                                 // PIXEL_GRABBER_RGB:sink_ready -> avalon_st_adapter_002:out_0_ready
	wire         avalon_st_adapter_002_out_0_startofpacket;                         // avalon_st_adapter_002:out_0_startofpacket -> PIXEL_GRABBER_RGB:sink_sop
	wire         avalon_st_adapter_002_out_0_endofpacket;                           // avalon_st_adapter_002:out_0_endofpacket -> PIXEL_GRABBER_RGB:sink_eop
	wire         dc_fifo_1_out_valid;                                               // dc_fifo_1:out_valid -> avalon_st_adapter_003:in_0_valid
	wire  [23:0] dc_fifo_1_out_data;                                                // dc_fifo_1:out_data -> avalon_st_adapter_003:in_0_data
	wire         dc_fifo_1_out_ready;                                               // avalon_st_adapter_003:in_0_ready -> dc_fifo_1:out_ready
	wire         dc_fifo_1_out_startofpacket;                                       // dc_fifo_1:out_startofpacket -> avalon_st_adapter_003:in_0_startofpacket
	wire         dc_fifo_1_out_endofpacket;                                         // dc_fifo_1:out_endofpacket -> avalon_st_adapter_003:in_0_endofpacket
	wire   [1:0] dc_fifo_1_out_empty;                                               // dc_fifo_1:out_empty -> avalon_st_adapter_003:in_0_empty
	wire         avalon_st_adapter_003_out_0_valid;                                 // avalon_st_adapter_003:out_0_valid -> data_format_adapter_0:in_valid
	wire  [23:0] avalon_st_adapter_003_out_0_data;                                  // avalon_st_adapter_003:out_0_data -> data_format_adapter_0:in_data
	wire         avalon_st_adapter_003_out_0_ready;                                 // data_format_adapter_0:in_ready -> avalon_st_adapter_003:out_0_ready
	wire         avalon_st_adapter_003_out_0_startofpacket;                         // avalon_st_adapter_003:out_0_startofpacket -> data_format_adapter_0:in_startofpacket
	wire         avalon_st_adapter_003_out_0_endofpacket;                           // avalon_st_adapter_003:out_0_endofpacket -> data_format_adapter_0:in_endofpacket
	wire   [1:0] avalon_st_adapter_003_out_0_empty;                                 // avalon_st_adapter_003:out_0_empty -> data_format_adapter_0:in_empty
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [COLOR_FILTER_0:reset_n, COM_COUNTER_0:reset_n, EDGE_BINS_0:reset_n, OBSTACLE_DIST_0:reset_n, PIXEL_BUFFER_0:reset_n, PIXEL_BUFFER_WB_0:reset_n, PIXEL_GRABBER_HSV:reset_n, PIXEL_GRABBER_RGB:reset_n, RGB_TO_HSV:reset_n, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, dc_fifo_0:out_reset_n, dc_fifo_1:in_reset_n, fir_0_0:main_reset, mm_interconnect_0:COLOR_FILTER_0_reset_reset_bridge_in_reset_reset]
	wire         nios2_gen2_debug_reset_request_reset;                              // nios2_gen2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [TERASIC_AUTO_FOCUS_0:reset_n, TERASIC_CAMERA_0:reset_n, alt_vip_itc_0:rst, alt_vip_vfb_0:reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, data_format_adapter_0:reset_n, dc_fifo_0:in_reset_n, dc_fifo_1:out_reset_n, mm_interconnect_0:TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:alt_vip_vfb_0_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [altpll_0:reset, altpll_2:reset, mm_interconnect_0:altpll_2_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                // rst_controller_003:reset_out -> [altpll_1:reset, i2c_opencores_camera:wb_rst_i, i2c_opencores_mipi:wb_rst_i, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, jtag_uart:rst_n, key:reset_n, led:reset_n, mipi_pwdn_n:reset_n, mipi_reset_n:reset_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, sw:reset_n, sysid_qsys:reset_n, uart_0:reset_n]
	wire         rst_controller_004_reset_out_reset;                                // rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, onchip_memory2_0:reset, pio_0:reset_n, rst_translator:in_reset, timer:reset_n, timer_0:reset_n]
	wire         rst_controller_004_reset_out_reset_req;                            // rst_controller_004:reset_req -> [nios2_gen2:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_005_reset_out_reset;                                // rst_controller_005:reset_out -> [mm_interconnect_0:timer_1_reset_reset_bridge_in_reset_reset, timer_1:reset_n]

	COLOR_FILTER color_filter_0 (
		.clk          (altpll_1_c0_clk),                                             //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                             //                   reset.reset_n
		.sink_data    (pixel_grabber_hsv_avalon_streaming_source_data),              //   avalon_streaming_sink.data
		.sink_eop     (pixel_grabber_hsv_avalon_streaming_source_endofpacket),       //                        .endofpacket
		.sink_ready   (pixel_grabber_hsv_avalon_streaming_source_ready),             //                        .ready
		.sink_sop     (pixel_grabber_hsv_avalon_streaming_source_startofpacket),     //                        .startofpacket
		.sink_valid   (pixel_grabber_hsv_avalon_streaming_source_valid),             //                        .valid
		.source_data  (color_filter_0_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (color_filter_0_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (color_filter_0_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (color_filter_0_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (color_filter_0_avalon_streaming_source_valid),                //                        .valid
		.s_chipselect (mm_interconnect_0_color_filter_0_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_color_filter_0_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_color_filter_0_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_color_filter_0_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_color_filter_0_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_color_filter_0_avalon_mm_slave_address)     //                        .address
	);

	COM_COUNTER_TOP #(
		.IMAGE_W (13'b0001010000000),
		.IMAGE_H (13'b0000111100000)
	) com_counter_0 (
		.clk          (altpll_1_c0_clk),                                            //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                            //                   reset.reset_n
		.sink_data    (fir_0_0_dout_data),                                          //   avalon_streaming_sink.data
		.sink_eop     (fir_0_0_dout_endofpacket),                                   //                        .endofpacket
		.sink_ready   (fir_0_0_dout_ready),                                         //                        .ready
		.sink_sop     (fir_0_0_dout_startofpacket),                                 //                        .startofpacket
		.sink_valid   (fir_0_0_dout_valid),                                         //                        .valid
		.source_data  (com_counter_0_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (com_counter_0_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (com_counter_0_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (com_counter_0_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (com_counter_0_avalon_streaming_source_valid),                //                        .valid
		.s_chipselect (mm_interconnect_0_com_counter_0_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_com_counter_0_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_com_counter_0_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_com_counter_0_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_com_counter_0_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_com_counter_0_avalon_mm_slave_address)     //                        .address
	);

	EDGE_BINS #(
		.IMAGE_W (13'b0001010000000),
		.IMAGE_H (13'b0000111100000)
	) edge_bins_0 (
		.clk          (altpll_1_c0_clk),                                          //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                          //                   reset.reset_n
		.source_data  (edge_bins_0_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (edge_bins_0_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (edge_bins_0_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (edge_bins_0_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (edge_bins_0_avalon_streaming_source_valid),                //                        .valid
		.sink_data    (com_counter_0_avalon_streaming_source_data),               //   avalon_streaming_sink.data
		.sink_valid   (com_counter_0_avalon_streaming_source_valid),              //                        .valid
		.sink_ready   (com_counter_0_avalon_streaming_source_ready),              //                        .ready
		.sink_sop     (com_counter_0_avalon_streaming_source_startofpacket),      //                        .startofpacket
		.sink_eop     (com_counter_0_avalon_streaming_source_endofpacket),        //                        .endofpacket
		.s_chipselect (mm_interconnect_0_edge_bins_0_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_edge_bins_0_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_edge_bins_0_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_edge_bins_0_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_edge_bins_0_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_edge_bins_0_avalon_mm_slave_address)     //                        .address
	);

	OBSTACLE_DIST #(
		.width  (640),
		.height (480)
	) obstacle_dist_0 (
		.clk          (altpll_1_c0_clk),                                              //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                              //                   reset.reset_n
		.s_chipselect (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_address),    //                        .address
		.sink_data    (edge_bins_0_avalon_streaming_source_data),                     //   avalon_streaming_sink.data
		.sink_eop     (edge_bins_0_avalon_streaming_source_endofpacket),              //                        .endofpacket
		.sink_ready   (edge_bins_0_avalon_streaming_source_ready),                    //                        .ready
		.sink_sop     (edge_bins_0_avalon_streaming_source_startofpacket),            //                        .startofpacket
		.sink_valid   (edge_bins_0_avalon_streaming_source_valid),                    //                        .valid
		.source_data  (obstacle_dist_0_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (obstacle_dist_0_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (obstacle_dist_0_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (obstacle_dist_0_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (obstacle_dist_0_avalon_streaming_source_valid)                 //                        .valid
	);

	PIXEL_BUFFER #(
		.width           (640),
		.height          (480),
		.sub_factor      (8),
		.clog_sub_factor (3)
	) pixel_buffer_0 (
		.clk          (altpll_1_c0_clk),                                             //                     clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.s_chipselect (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_chipselect), //           avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_read),       //                          .read
		.s_write      (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_write),      //                          .write
		.s_readdata   (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_readdata),   //                          .readdata
		.s_writedata  (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_writedata),  //                          .writedata
		.s_address    (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_address),    //                          .address
		.sink_data    (pixel_grabber_rgb_avalon_streaming_source_data),              //     avalon_streaming_sink.data
		.sink_eop     (pixel_grabber_rgb_avalon_streaming_source_endofpacket),       //                          .endofpacket
		.sink_ready   (pixel_grabber_rgb_avalon_streaming_source_ready),             //                          .ready
		.sink_sop     (pixel_grabber_rgb_avalon_streaming_source_startofpacket),     //                          .startofpacket
		.sink_valid   (pixel_grabber_rgb_avalon_streaming_source_valid),             //                          .valid
		.source_data  (pixel_buffer_0_avalon_streaming_source_1_data),               // avalon_streaming_source_1.data
		.source_eop   (pixel_buffer_0_avalon_streaming_source_1_endofpacket),        //                          .endofpacket
		.source_ready (pixel_buffer_0_avalon_streaming_source_1_ready),              //                          .ready
		.source_sop   (pixel_buffer_0_avalon_streaming_source_1_startofpacket),      //                          .startofpacket
		.source_valid (pixel_buffer_0_avalon_streaming_source_1_valid)               //                          .valid
	);

	PIXEL_BUFFER_WB #(
		.width           (640),
		.height          (480),
		.sub_factor      (32),
		.clog_sub_factor (5)
	) pixel_buffer_wb_0 (
		.clk          (altpll_1_c0_clk),                                                //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                                //                   reset.reset_n
		.s_chipselect (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_address),    //                        .address
		.sink_data    (pixel_buffer_0_avalon_streaming_source_1_data),                  //   avalon_streaming_sink.data
		.sink_eop     (pixel_buffer_0_avalon_streaming_source_1_endofpacket),           //                        .endofpacket
		.sink_ready   (pixel_buffer_0_avalon_streaming_source_1_ready),                 //                        .ready
		.sink_sop     (pixel_buffer_0_avalon_streaming_source_1_startofpacket),         //                        .startofpacket
		.sink_valid   (pixel_buffer_0_avalon_streaming_source_1_valid),                 //                        .valid
		.source_data  (pixel_buffer_wb_0_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (pixel_buffer_wb_0_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (pixel_buffer_wb_0_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (pixel_buffer_wb_0_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (pixel_buffer_wb_0_avalon_streaming_source_valid)                 //                        .valid
	);

	PIXEL_GRABBER #(
		.width  (640),
		.height (480)
	) pixel_grabber_hsv (
		.clk          (altpll_1_c0_clk),                                                //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                                //                   reset.reset_n
		.sink_data    (rgb_to_hsv_avalon_streaming_source_data),                        //   avalon_streaming_sink.data
		.sink_eop     (rgb_to_hsv_avalon_streaming_source_endofpacket),                 //                        .endofpacket
		.sink_ready   (rgb_to_hsv_avalon_streaming_source_ready),                       //                        .ready
		.sink_sop     (rgb_to_hsv_avalon_streaming_source_startofpacket),               //                        .startofpacket
		.sink_valid   (rgb_to_hsv_avalon_streaming_source_valid),                       //                        .valid
		.source_data  (pixel_grabber_hsv_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (pixel_grabber_hsv_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (pixel_grabber_hsv_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (pixel_grabber_hsv_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (pixel_grabber_hsv_avalon_streaming_source_valid),                //                        .valid
		.s_chipselect (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_address)     //                        .address
	);

	PIXEL_GRABBER #(
		.width  (640),
		.height (480)
	) pixel_grabber_rgb (
		.clk          (altpll_1_c0_clk),                                                //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                                //                   reset.reset_n
		.sink_data    (avalon_st_adapter_002_out_0_data),                               //   avalon_streaming_sink.data
		.sink_eop     (avalon_st_adapter_002_out_0_endofpacket),                        //                        .endofpacket
		.sink_ready   (avalon_st_adapter_002_out_0_ready),                              //                        .ready
		.sink_sop     (avalon_st_adapter_002_out_0_startofpacket),                      //                        .startofpacket
		.sink_valid   (avalon_st_adapter_002_out_0_valid),                              //                        .valid
		.source_data  (pixel_grabber_rgb_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (pixel_grabber_rgb_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (pixel_grabber_rgb_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (pixel_grabber_rgb_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (pixel_grabber_rgb_avalon_streaming_source_valid),                //                        .valid
		.s_chipselect (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_address)     //                        .address
	);

	RGB_TO_HSV_PIPELINED_TOP rgb_to_hsv (
		.clk          (altpll_1_c0_clk),                                         //                   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                         //                   reset.reset_n
		.sink_data    (pixel_buffer_wb_0_avalon_streaming_source_data),          //   avalon_streaming_sink.data
		.sink_eop     (pixel_buffer_wb_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.sink_ready   (pixel_buffer_wb_0_avalon_streaming_source_ready),         //                        .ready
		.sink_sop     (pixel_buffer_wb_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.sink_valid   (pixel_buffer_wb_0_avalon_streaming_source_valid),         //                        .valid
		.source_data  (rgb_to_hsv_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.source_eop   (rgb_to_hsv_avalon_streaming_source_endofpacket),          //                        .endofpacket
		.source_ready (rgb_to_hsv_avalon_streaming_source_ready),                //                        .ready
		.source_sop   (rgb_to_hsv_avalon_streaming_source_startofpacket),        //                        .startofpacket
		.source_valid (rgb_to_hsv_avalon_streaming_source_valid),                //                        .valid
		.s_chipselect (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_chipselect), //         avalon_mm_slave.chipselect
		.s_read       (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_read),       //                        .read
		.s_write      (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_write),      //                        .write
		.s_readdata   (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_readdata),   //                        .readdata
		.s_writedata  (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_writedata),  //                        .writedata
		.s_address    (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_address)     //                        .address
	);

	TERASIC_AUTO_FOCUS #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_auto_focus_0 (
		.clk          (altpll_0_c2_clk),                                           //   clock.clk
		.reset_n      (~rst_controller_001_reset_out_reset),                       //   reset.reset_n
		.s_chipselect (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect), // mm_ctrl.chipselect
		.s_read       (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read),       //        .read
		.s_write      (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write),      //        .write
		.s_readdata   (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata),   //        .readdata
		.s_writedata  (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata),  //        .writedata
		.s_address    (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address),    //        .address
		.sink_data    (alt_vip_vfb_0_dout_data),                                   //     din.data
		.sink_valid   (alt_vip_vfb_0_dout_valid),                                  //        .valid
		.sink_ready   (alt_vip_vfb_0_dout_ready),                                  //        .ready
		.sink_sop     (alt_vip_vfb_0_dout_startofpacket),                          //        .startofpacket
		.sink_eop     (alt_vip_vfb_0_dout_endofpacket),                            //        .endofpacket
		.source_data  (terasic_auto_focus_0_dout_data),                            //    dout.data
		.source_valid (terasic_auto_focus_0_dout_valid),                           //        .valid
		.source_ready (terasic_auto_focus_0_dout_ready),                           //        .ready
		.source_sop   (terasic_auto_focus_0_dout_startofpacket),                   //        .startofpacket
		.source_eop   (terasic_auto_focus_0_dout_endofpacket),                     //        .endofpacket
		.vcm_i2c_sda  (terasic_auto_focus_0_conduit_vcm_i2c_sda),                  // Conduit.vcm_i2c_sda
		.clk50        (terasic_auto_focus_0_conduit_clk50),                        //        .clk50
		.vcm_i2c_scl  (terasic_auto_focus_0_conduit_vcm_i2c_scl)                   //        .vcm_i2c_scl
	);

	TERASIC_CAMERA #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_camera_0 (
		.clk           (altpll_0_c2_clk),                                        //             clock_reset.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //       clock_reset_reset.reset_n
		.CAMERA_D      (terasic_camera_0_conduit_end_D),                         //             conduit_end.export
		.CAMERA_FVAL   (terasic_camera_0_conduit_end_FVAL),                      //                        .export
		.CAMERA_LVAL   (terasic_camera_0_conduit_end_LVAL),                      //                        .export
		.CAMERA_PIXCLK (terasic_camera_0_conduit_end_PIXCLK),                    //                        .export
		.st_data       (terasic_camera_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.st_sop        (terasic_camera_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.st_eop        (terasic_camera_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.st_ready      (terasic_camera_0_avalon_streaming_source_ready),         //                        .ready
		.st_valid      (terasic_camera_0_avalon_streaming_source_valid)          //                        .valid
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (640),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (640),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (639),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (96),
		.H_FRONT_PORCH                 (16),
		.H_BACK_PORCH                  (48),
		.V_SYNC_LENGTH                 (2),
		.V_FRONT_PORCH                 (10),
		.V_BACK_PORCH                  (33),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (altpll_0_c2_clk),                           //       is_clk_rst.clk
		.rst           (rst_controller_001_reset_out_reset),        // is_clk_rst_reset.reset
		.is_data       (data_format_adapter_0_out_data),            //              din.data
		.is_valid      (data_format_adapter_0_out_valid),           //                 .valid
		.is_ready      (data_format_adapter_0_out_ready),           //                 .ready
		.is_sop        (data_format_adapter_0_out_startofpacket),   //                 .startofpacket
		.is_eop        (data_format_adapter_0_out_endofpacket),     //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	Qsys_alt_vip_vfb_0 alt_vip_vfb_0 (
		.clock                        (altpll_0_c2_clk),                                        //        clock.clk
		.reset                        (rst_controller_001_reset_out_reset),                     //        reset.reset
		.din_ready                    (terasic_camera_0_avalon_streaming_source_ready),         //          din.ready
		.din_valid                    (terasic_camera_0_avalon_streaming_source_valid),         //             .valid
		.din_data                     (terasic_camera_0_avalon_streaming_source_data),          //             .data
		.din_startofpacket            (terasic_camera_0_avalon_streaming_source_startofpacket), //             .startofpacket
		.din_endofpacket              (terasic_camera_0_avalon_streaming_source_endofpacket),   //             .endofpacket
		.dout_ready                   (alt_vip_vfb_0_dout_ready),                               //         dout.ready
		.dout_valid                   (alt_vip_vfb_0_dout_valid),                               //             .valid
		.dout_data                    (alt_vip_vfb_0_dout_data),                                //             .data
		.dout_startofpacket           (alt_vip_vfb_0_dout_startofpacket),                       //             .startofpacket
		.dout_endofpacket             (alt_vip_vfb_0_dout_endofpacket),                         //             .endofpacket
		.read_master_av_address       (alt_vip_vfb_0_read_master_address),                      //  read_master.address
		.read_master_av_read          (alt_vip_vfb_0_read_master_read),                         //             .read
		.read_master_av_waitrequest   (alt_vip_vfb_0_read_master_waitrequest),                  //             .waitrequest
		.read_master_av_readdatavalid (alt_vip_vfb_0_read_master_readdatavalid),                //             .readdatavalid
		.read_master_av_readdata      (alt_vip_vfb_0_read_master_readdata),                     //             .readdata
		.read_master_av_burstcount    (alt_vip_vfb_0_read_master_burstcount),                   //             .burstcount
		.write_master_av_address      (alt_vip_vfb_0_write_master_address),                     // write_master.address
		.write_master_av_write        (alt_vip_vfb_0_write_master_write),                       //             .write
		.write_master_av_writedata    (alt_vip_vfb_0_write_master_writedata),                   //             .writedata
		.write_master_av_waitrequest  (alt_vip_vfb_0_write_master_waitrequest),                 //             .waitrequest
		.write_master_av_burstcount   (alt_vip_vfb_0_write_master_burstcount)                   //             .burstcount
	);

	Qsys_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (),                                               //                    c0.clk
		.c1                 (clk_sdram_clk),                                  //                    c1.clk
		.c2                 (altpll_0_c2_clk),                                //                    c2.clk
		.c3                 (clk_vga_clk),                                    //                    c3.clk
		.c4                 (d8m_xclkin_clk),                                 //                    c4.clk
		.areset             (altpll_0_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_0_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	Qsys_altpll_1 altpll_1 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_003_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_1_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_1_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_1_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_1_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_1_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_1_c0_clk),                                //                    c0.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c1                 (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	Qsys_altpll_2 altpll_2 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_2_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_2_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_2_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_2_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_2_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_2_c0_clk),                                //                    c0.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c1                 (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	Qsys_data_format_adapter_0 data_format_adapter_0 (
		.clk               (altpll_0_c2_clk),                           //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset),       // reset.reset_n
		.in_data           (avalon_st_adapter_003_out_0_data),          //    in.data
		.in_valid          (avalon_st_adapter_003_out_0_valid),         //      .valid
		.in_ready          (avalon_st_adapter_003_out_0_ready),         //      .ready
		.in_startofpacket  (avalon_st_adapter_003_out_0_startofpacket), //      .startofpacket
		.in_endofpacket    (avalon_st_adapter_003_out_0_endofpacket),   //      .endofpacket
		.in_empty          (avalon_st_adapter_003_out_0_empty),         //      .empty
		.out_data          (data_format_adapter_0_out_data),            //   out.data
		.out_valid         (data_format_adapter_0_out_valid),           //      .valid
		.out_ready         (data_format_adapter_0_out_ready),           //      .ready
		.out_startofpacket (data_format_adapter_0_out_startofpacket),   //      .startofpacket
		.out_endofpacket   (data_format_adapter_0_out_endofpacket)      //      .endofpacket
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (3),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (128),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dc_fifo_0 (
		.in_clk            (altpll_0_c2_clk),                           //        in_clk.clk
		.in_reset_n        (~rst_controller_001_reset_out_reset),       //  in_clk_reset.reset_n
		.out_clk           (altpll_1_c0_clk),                           //       out_clk.clk
		.out_reset_n       (~rst_controller_reset_out_reset),           // out_clk_reset.reset_n
		.in_data           (avalon_st_adapter_001_out_0_data),          //            in.data
		.in_valid          (avalon_st_adapter_001_out_0_valid),         //              .valid
		.in_ready          (avalon_st_adapter_001_out_0_ready),         //              .ready
		.in_startofpacket  (avalon_st_adapter_001_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_001_out_0_endofpacket),   //              .endofpacket
		.in_empty          (avalon_st_adapter_001_out_0_empty),         //              .empty
		.out_data          (dc_fifo_0_out_data),                        //           out.data
		.out_valid         (dc_fifo_0_out_valid),                       //              .valid
		.out_ready         (dc_fifo_0_out_ready),                       //              .ready
		.out_startofpacket (dc_fifo_0_out_startofpacket),               //              .startofpacket
		.out_endofpacket   (dc_fifo_0_out_endofpacket),                 //              .endofpacket
		.out_empty         (dc_fifo_0_out_empty),                       //              .empty
		.in_csr_address    (1'b0),                                      //   (terminated)
		.in_csr_read       (1'b0),                                      //   (terminated)
		.in_csr_write      (1'b0),                                      //   (terminated)
		.in_csr_readdata   (),                                          //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),      //   (terminated)
		.out_csr_address   (1'b0),                                      //   (terminated)
		.out_csr_read      (1'b0),                                      //   (terminated)
		.out_csr_write     (1'b0),                                      //   (terminated)
		.out_csr_readdata  (),                                          //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000),      //   (terminated)
		.in_error          (1'b0),                                      //   (terminated)
		.out_error         (),                                          //   (terminated)
		.in_channel        (1'b0),                                      //   (terminated)
		.out_channel       (),                                          //   (terminated)
		.space_avail_data  ()                                           //   (terminated)
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (3),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (128),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dc_fifo_1 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),       //  in_clk_reset.reset_n
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),   // out_clk_reset.reset_n
		.in_data           (avalon_st_adapter_out_0_data),          //            in.data
		.in_valid          (avalon_st_adapter_out_0_valid),         //              .valid
		.in_ready          (avalon_st_adapter_out_0_ready),         //              .ready
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //              .endofpacket
		.in_empty          (avalon_st_adapter_out_0_empty),         //              .empty
		.out_data          (dc_fifo_1_out_data),                    //           out.data
		.out_valid         (dc_fifo_1_out_valid),                   //              .valid
		.out_ready         (dc_fifo_1_out_ready),                   //              .ready
		.out_startofpacket (dc_fifo_1_out_startofpacket),           //              .startofpacket
		.out_endofpacket   (dc_fifo_1_out_endofpacket),             //              .endofpacket
		.out_empty         (dc_fifo_1_out_empty),                   //              .empty
		.in_csr_address    (1'b0),                                  //   (terminated)
		.in_csr_read       (1'b0),                                  //   (terminated)
		.in_csr_write      (1'b0),                                  //   (terminated)
		.in_csr_readdata   (),                                      //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),  //   (terminated)
		.out_csr_address   (1'b0),                                  //   (terminated)
		.out_csr_read      (1'b0),                                  //   (terminated)
		.out_csr_write     (1'b0),                                  //   (terminated)
		.out_csr_readdata  (),                                      //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000),  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_error         (),                                      //   (terminated)
		.in_channel        (1'b0),                                  //   (terminated)
		.out_channel       (),                                      //   (terminated)
		.space_avail_data  ()                                       //   (terminated)
	);

	Qsys_fir_0_0 fir_0_0 (
		.main_clock            (altpll_1_c0_clk),                                      // main_clock.clk
		.main_reset            (rst_controller_reset_out_reset),                       // main_reset.reset
		.din_data              (color_filter_0_avalon_streaming_source_data),          //        din.data
		.din_valid             (color_filter_0_avalon_streaming_source_valid),         //           .valid
		.din_startofpacket     (color_filter_0_avalon_streaming_source_startofpacket), //           .startofpacket
		.din_endofpacket       (color_filter_0_avalon_streaming_source_endofpacket),   //           .endofpacket
		.din_ready             (color_filter_0_avalon_streaming_source_ready),         //           .ready
		.dout_data             (fir_0_0_dout_data),                                    //       dout.data
		.dout_valid            (fir_0_0_dout_valid),                                   //           .valid
		.dout_startofpacket    (fir_0_0_dout_startofpacket),                           //           .startofpacket
		.dout_endofpacket      (fir_0_0_dout_endofpacket),                             //           .endofpacket
		.dout_ready            (fir_0_0_dout_ready),                                   //           .ready
		.control_address       (mm_interconnect_0_fir_0_0_control_address),            //    control.address
		.control_byteenable    (mm_interconnect_0_fir_0_0_control_byteenable),         //           .byteenable
		.control_write         (mm_interconnect_0_fir_0_0_control_write),              //           .write
		.control_writedata     (mm_interconnect_0_fir_0_0_control_writedata),          //           .writedata
		.control_read          (mm_interconnect_0_fir_0_0_control_read),               //           .read
		.control_readdata      (mm_interconnect_0_fir_0_0_control_readdata),           //           .readdata
		.control_readdatavalid (mm_interconnect_0_fir_0_0_control_readdatavalid),      //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_fir_0_0_control_waitrequest)         //           .waitrequest
	);

	i2c_opencores i2c_opencores_camera (
		.wb_clk_i   (clk_clk),                                                           //            clock.clk
		.wb_rst_i   (rst_controller_003_reset_out_reset),                                //      clock_reset.reset
		.scl_pad_io (i2c_opencores_camera_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_camera_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_001_receiver_irq)                                  // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_mipi (
		.wb_clk_i   (clk_clk),                                                         //            clock.clk
		.wb_rst_i   (rst_controller_003_reset_out_reset),                              //      clock_reset.reset
		.scl_pad_io (i2c_opencores_mipi_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_mipi_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_receiver_irq)                                    // interrupt_sender.irq
	);

	Qsys_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_002_receiver_irq)                          //               irq.irq
	);

	Qsys_key key (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	Qsys_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	Qsys_mipi_pwdn_n mipi_pwdn_n (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mipi_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_pwdn_n_external_connection_export)       // external_connection.export
	);

	Qsys_mipi_pwdn_n mipi_reset_n (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_external_connection_export)       // external_connection.export
	);

	Qsys_nios2_gen2 nios2_gen2 (
		.clk                                 (altpll_2_c0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_004_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_004_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	Qsys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_2_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_004_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	Qsys_pio_0 pio_0 (
		.clk        (altpll_2_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.in_port    (switch_export),                         // external_connection.export
		.irq        (irq_mapper_receiver6_irq)               //                 irq.irq
	);

	Qsys_sdram sdram (
		.clk            (altpll_0_c2_clk),                          //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Qsys_sw sw (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata),    //                    .readdata
		.in_port  (sw_external_connection_export)        // external_connection.export
	);

	Qsys_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	Qsys_timer timer (
		.clk        (altpll_2_c0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
	);

	Qsys_timer_0 timer_0 (
		.clk        (altpll_2_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	Qsys_timer_0 timer_1 (
		.clk        (altpll_2_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver7_irq)                 //   irq.irq
	);

	Qsys_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_003_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_rx_tx_rxd),                          // external_connection.export
		.txd           (uart_0_rx_tx_txd),                          //                    .export
		.irq           (irq_synchronizer_003_receiver_irq)          //                 irq.irq
	);

	Qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c2_clk                                            (altpll_0_c2_clk),                                                    //                                          altpll_0_c2.clk
		.altpll_1_c0_clk                                            (altpll_1_c0_clk),                                                    //                                          altpll_1_c0.clk
		.altpll_2_c0_clk                                            (altpll_2_c0_clk),                                                    //                                          altpll_2_c0.clk
		.clk_50_clk_clk                                             (clk_clk),                                                            //                                           clk_50_clk.clk
		.altpll_2_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                 // altpll_2_inclk_interface_reset_reset_bridge_in_reset.reset
		.COLOR_FILTER_0_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                     //           COLOR_FILTER_0_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset                (rst_controller_003_reset_out_reset),                                 //                jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset               (rst_controller_004_reset_out_reset),                                 //               nios2_gen2_reset_reset_bridge_in_reset.reset
		.TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                 //     TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset.reset
		.timer_1_reset_reset_bridge_in_reset_reset                  (rst_controller_005_reset_out_reset),                                 //                  timer_1_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                             (nios2_gen2_data_master_address),                                     //                               nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                         (nios2_gen2_data_master_waitrequest),                                 //                                                     .waitrequest
		.nios2_gen2_data_master_byteenable                          (nios2_gen2_data_master_byteenable),                                  //                                                     .byteenable
		.nios2_gen2_data_master_read                                (nios2_gen2_data_master_read),                                        //                                                     .read
		.nios2_gen2_data_master_readdata                            (nios2_gen2_data_master_readdata),                                    //                                                     .readdata
		.nios2_gen2_data_master_readdatavalid                       (nios2_gen2_data_master_readdatavalid),                               //                                                     .readdatavalid
		.nios2_gen2_data_master_write                               (nios2_gen2_data_master_write),                                       //                                                     .write
		.nios2_gen2_data_master_writedata                           (nios2_gen2_data_master_writedata),                                   //                                                     .writedata
		.nios2_gen2_data_master_debugaccess                         (nios2_gen2_data_master_debugaccess),                                 //                                                     .debugaccess
		.nios2_gen2_instruction_master_address                      (nios2_gen2_instruction_master_address),                              //                        nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                  (nios2_gen2_instruction_master_waitrequest),                          //                                                     .waitrequest
		.nios2_gen2_instruction_master_read                         (nios2_gen2_instruction_master_read),                                 //                                                     .read
		.nios2_gen2_instruction_master_readdata                     (nios2_gen2_instruction_master_readdata),                             //                                                     .readdata
		.nios2_gen2_instruction_master_readdatavalid                (nios2_gen2_instruction_master_readdatavalid),                        //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                       //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                         //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                          //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                      //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                     //                                                     .writedata
		.altpll_1_pll_slave_address                                 (mm_interconnect_0_altpll_1_pll_slave_address),                       //                                   altpll_1_pll_slave.address
		.altpll_1_pll_slave_write                                   (mm_interconnect_0_altpll_1_pll_slave_write),                         //                                                     .write
		.altpll_1_pll_slave_read                                    (mm_interconnect_0_altpll_1_pll_slave_read),                          //                                                     .read
		.altpll_1_pll_slave_readdata                                (mm_interconnect_0_altpll_1_pll_slave_readdata),                      //                                                     .readdata
		.altpll_1_pll_slave_writedata                               (mm_interconnect_0_altpll_1_pll_slave_writedata),                     //                                                     .writedata
		.altpll_2_pll_slave_address                                 (mm_interconnect_0_altpll_2_pll_slave_address),                       //                                   altpll_2_pll_slave.address
		.altpll_2_pll_slave_write                                   (mm_interconnect_0_altpll_2_pll_slave_write),                         //                                                     .write
		.altpll_2_pll_slave_read                                    (mm_interconnect_0_altpll_2_pll_slave_read),                          //                                                     .read
		.altpll_2_pll_slave_readdata                                (mm_interconnect_0_altpll_2_pll_slave_readdata),                      //                                                     .readdata
		.altpll_2_pll_slave_writedata                               (mm_interconnect_0_altpll_2_pll_slave_writedata),                     //                                                     .writedata
		.COLOR_FILTER_0_avalon_mm_slave_address                     (mm_interconnect_0_color_filter_0_avalon_mm_slave_address),           //                       COLOR_FILTER_0_avalon_mm_slave.address
		.COLOR_FILTER_0_avalon_mm_slave_write                       (mm_interconnect_0_color_filter_0_avalon_mm_slave_write),             //                                                     .write
		.COLOR_FILTER_0_avalon_mm_slave_read                        (mm_interconnect_0_color_filter_0_avalon_mm_slave_read),              //                                                     .read
		.COLOR_FILTER_0_avalon_mm_slave_readdata                    (mm_interconnect_0_color_filter_0_avalon_mm_slave_readdata),          //                                                     .readdata
		.COLOR_FILTER_0_avalon_mm_slave_writedata                   (mm_interconnect_0_color_filter_0_avalon_mm_slave_writedata),         //                                                     .writedata
		.COLOR_FILTER_0_avalon_mm_slave_chipselect                  (mm_interconnect_0_color_filter_0_avalon_mm_slave_chipselect),        //                                                     .chipselect
		.COM_COUNTER_0_avalon_mm_slave_address                      (mm_interconnect_0_com_counter_0_avalon_mm_slave_address),            //                        COM_COUNTER_0_avalon_mm_slave.address
		.COM_COUNTER_0_avalon_mm_slave_write                        (mm_interconnect_0_com_counter_0_avalon_mm_slave_write),              //                                                     .write
		.COM_COUNTER_0_avalon_mm_slave_read                         (mm_interconnect_0_com_counter_0_avalon_mm_slave_read),               //                                                     .read
		.COM_COUNTER_0_avalon_mm_slave_readdata                     (mm_interconnect_0_com_counter_0_avalon_mm_slave_readdata),           //                                                     .readdata
		.COM_COUNTER_0_avalon_mm_slave_writedata                    (mm_interconnect_0_com_counter_0_avalon_mm_slave_writedata),          //                                                     .writedata
		.COM_COUNTER_0_avalon_mm_slave_chipselect                   (mm_interconnect_0_com_counter_0_avalon_mm_slave_chipselect),         //                                                     .chipselect
		.EDGE_BINS_0_avalon_mm_slave_address                        (mm_interconnect_0_edge_bins_0_avalon_mm_slave_address),              //                          EDGE_BINS_0_avalon_mm_slave.address
		.EDGE_BINS_0_avalon_mm_slave_write                          (mm_interconnect_0_edge_bins_0_avalon_mm_slave_write),                //                                                     .write
		.EDGE_BINS_0_avalon_mm_slave_read                           (mm_interconnect_0_edge_bins_0_avalon_mm_slave_read),                 //                                                     .read
		.EDGE_BINS_0_avalon_mm_slave_readdata                       (mm_interconnect_0_edge_bins_0_avalon_mm_slave_readdata),             //                                                     .readdata
		.EDGE_BINS_0_avalon_mm_slave_writedata                      (mm_interconnect_0_edge_bins_0_avalon_mm_slave_writedata),            //                                                     .writedata
		.EDGE_BINS_0_avalon_mm_slave_chipselect                     (mm_interconnect_0_edge_bins_0_avalon_mm_slave_chipselect),           //                                                     .chipselect
		.fir_0_0_control_address                                    (mm_interconnect_0_fir_0_0_control_address),                          //                                      fir_0_0_control.address
		.fir_0_0_control_write                                      (mm_interconnect_0_fir_0_0_control_write),                            //                                                     .write
		.fir_0_0_control_read                                       (mm_interconnect_0_fir_0_0_control_read),                             //                                                     .read
		.fir_0_0_control_readdata                                   (mm_interconnect_0_fir_0_0_control_readdata),                         //                                                     .readdata
		.fir_0_0_control_writedata                                  (mm_interconnect_0_fir_0_0_control_writedata),                        //                                                     .writedata
		.fir_0_0_control_byteenable                                 (mm_interconnect_0_fir_0_0_control_byteenable),                       //                                                     .byteenable
		.fir_0_0_control_readdatavalid                              (mm_interconnect_0_fir_0_0_control_readdatavalid),                    //                                                     .readdatavalid
		.fir_0_0_control_waitrequest                                (mm_interconnect_0_fir_0_0_control_waitrequest),                      //                                                     .waitrequest
		.i2c_opencores_camera_avalon_slave_0_address                (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address),      //                  i2c_opencores_camera_avalon_slave_0.address
		.i2c_opencores_camera_avalon_slave_0_write                  (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write),        //                                                     .write
		.i2c_opencores_camera_avalon_slave_0_readdata               (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata),     //                                                     .readdata
		.i2c_opencores_camera_avalon_slave_0_writedata              (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata),    //                                                     .writedata
		.i2c_opencores_camera_avalon_slave_0_waitrequest            (~mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest), //                                                     .waitrequest
		.i2c_opencores_camera_avalon_slave_0_chipselect             (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect),   //                                                     .chipselect
		.i2c_opencores_mipi_avalon_slave_0_address                  (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address),        //                    i2c_opencores_mipi_avalon_slave_0.address
		.i2c_opencores_mipi_avalon_slave_0_write                    (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write),          //                                                     .write
		.i2c_opencores_mipi_avalon_slave_0_readdata                 (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata),       //                                                     .readdata
		.i2c_opencores_mipi_avalon_slave_0_writedata                (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata),      //                                                     .writedata
		.i2c_opencores_mipi_avalon_slave_0_waitrequest              (~mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest),   //                                                     .waitrequest
		.i2c_opencores_mipi_avalon_slave_0_chipselect               (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect),     //                                                     .chipselect
		.jtag_uart_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                                     .chipselect
		.key_s1_address                                             (mm_interconnect_0_key_s1_address),                                   //                                               key_s1.address
		.key_s1_readdata                                            (mm_interconnect_0_key_s1_readdata),                                  //                                                     .readdata
		.led_s1_address                                             (mm_interconnect_0_led_s1_address),                                   //                                               led_s1.address
		.led_s1_write                                               (mm_interconnect_0_led_s1_write),                                     //                                                     .write
		.led_s1_readdata                                            (mm_interconnect_0_led_s1_readdata),                                  //                                                     .readdata
		.led_s1_writedata                                           (mm_interconnect_0_led_s1_writedata),                                 //                                                     .writedata
		.led_s1_chipselect                                          (mm_interconnect_0_led_s1_chipselect),                                //                                                     .chipselect
		.mipi_pwdn_n_s1_address                                     (mm_interconnect_0_mipi_pwdn_n_s1_address),                           //                                       mipi_pwdn_n_s1.address
		.mipi_pwdn_n_s1_write                                       (mm_interconnect_0_mipi_pwdn_n_s1_write),                             //                                                     .write
		.mipi_pwdn_n_s1_readdata                                    (mm_interconnect_0_mipi_pwdn_n_s1_readdata),                          //                                                     .readdata
		.mipi_pwdn_n_s1_writedata                                   (mm_interconnect_0_mipi_pwdn_n_s1_writedata),                         //                                                     .writedata
		.mipi_pwdn_n_s1_chipselect                                  (mm_interconnect_0_mipi_pwdn_n_s1_chipselect),                        //                                                     .chipselect
		.mipi_reset_n_s1_address                                    (mm_interconnect_0_mipi_reset_n_s1_address),                          //                                      mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                                      (mm_interconnect_0_mipi_reset_n_s1_write),                            //                                                     .write
		.mipi_reset_n_s1_readdata                                   (mm_interconnect_0_mipi_reset_n_s1_readdata),                         //                                                     .readdata
		.mipi_reset_n_s1_writedata                                  (mm_interconnect_0_mipi_reset_n_s1_writedata),                        //                                                     .writedata
		.mipi_reset_n_s1_chipselect                                 (mm_interconnect_0_mipi_reset_n_s1_chipselect),                       //                                                     .chipselect
		.nios2_gen2_debug_mem_slave_address                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),               //                           nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                           (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),                 //                                                     .write
		.nios2_gen2_debug_mem_slave_read                            (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),                  //                                                     .read
		.nios2_gen2_debug_mem_slave_readdata                        (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),              //                                                     .readdata
		.nios2_gen2_debug_mem_slave_writedata                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),             //                                                     .writedata
		.nios2_gen2_debug_mem_slave_byteenable                      (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),            //                                                     .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),           //                                                     .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),           //                                                     .debugaccess
		.OBSTACLE_DIST_0_avalon_mm_slave_address                    (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_address),          //                      OBSTACLE_DIST_0_avalon_mm_slave.address
		.OBSTACLE_DIST_0_avalon_mm_slave_write                      (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_write),            //                                                     .write
		.OBSTACLE_DIST_0_avalon_mm_slave_read                       (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_read),             //                                                     .read
		.OBSTACLE_DIST_0_avalon_mm_slave_readdata                   (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_readdata),         //                                                     .readdata
		.OBSTACLE_DIST_0_avalon_mm_slave_writedata                  (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_writedata),        //                                                     .writedata
		.OBSTACLE_DIST_0_avalon_mm_slave_chipselect                 (mm_interconnect_0_obstacle_dist_0_avalon_mm_slave_chipselect),       //                                                     .chipselect
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                      //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                        //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                     //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),                    //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                   //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                   //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                        //                                                     .clken
		.pio_0_s1_address                                           (mm_interconnect_0_pio_0_s1_address),                                 //                                             pio_0_s1.address
		.pio_0_s1_write                                             (mm_interconnect_0_pio_0_s1_write),                                   //                                                     .write
		.pio_0_s1_readdata                                          (mm_interconnect_0_pio_0_s1_readdata),                                //                                                     .readdata
		.pio_0_s1_writedata                                         (mm_interconnect_0_pio_0_s1_writedata),                               //                                                     .writedata
		.pio_0_s1_chipselect                                        (mm_interconnect_0_pio_0_s1_chipselect),                              //                                                     .chipselect
		.PIXEL_BUFFER_0_avalon_mm_slave_address                     (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_address),           //                       PIXEL_BUFFER_0_avalon_mm_slave.address
		.PIXEL_BUFFER_0_avalon_mm_slave_write                       (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_write),             //                                                     .write
		.PIXEL_BUFFER_0_avalon_mm_slave_read                        (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_read),              //                                                     .read
		.PIXEL_BUFFER_0_avalon_mm_slave_readdata                    (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_readdata),          //                                                     .readdata
		.PIXEL_BUFFER_0_avalon_mm_slave_writedata                   (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_writedata),         //                                                     .writedata
		.PIXEL_BUFFER_0_avalon_mm_slave_chipselect                  (mm_interconnect_0_pixel_buffer_0_avalon_mm_slave_chipselect),        //                                                     .chipselect
		.PIXEL_BUFFER_WB_0_avalon_mm_slave_address                  (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_address),        //                    PIXEL_BUFFER_WB_0_avalon_mm_slave.address
		.PIXEL_BUFFER_WB_0_avalon_mm_slave_write                    (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_write),          //                                                     .write
		.PIXEL_BUFFER_WB_0_avalon_mm_slave_read                     (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_read),           //                                                     .read
		.PIXEL_BUFFER_WB_0_avalon_mm_slave_readdata                 (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_readdata),       //                                                     .readdata
		.PIXEL_BUFFER_WB_0_avalon_mm_slave_writedata                (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_writedata),      //                                                     .writedata
		.PIXEL_BUFFER_WB_0_avalon_mm_slave_chipselect               (mm_interconnect_0_pixel_buffer_wb_0_avalon_mm_slave_chipselect),     //                                                     .chipselect
		.PIXEL_GRABBER_HSV_avalon_mm_slave_address                  (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_address),        //                    PIXEL_GRABBER_HSV_avalon_mm_slave.address
		.PIXEL_GRABBER_HSV_avalon_mm_slave_write                    (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_write),          //                                                     .write
		.PIXEL_GRABBER_HSV_avalon_mm_slave_read                     (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_read),           //                                                     .read
		.PIXEL_GRABBER_HSV_avalon_mm_slave_readdata                 (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_readdata),       //                                                     .readdata
		.PIXEL_GRABBER_HSV_avalon_mm_slave_writedata                (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_writedata),      //                                                     .writedata
		.PIXEL_GRABBER_HSV_avalon_mm_slave_chipselect               (mm_interconnect_0_pixel_grabber_hsv_avalon_mm_slave_chipselect),     //                                                     .chipselect
		.PIXEL_GRABBER_RGB_avalon_mm_slave_address                  (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_address),        //                    PIXEL_GRABBER_RGB_avalon_mm_slave.address
		.PIXEL_GRABBER_RGB_avalon_mm_slave_write                    (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_write),          //                                                     .write
		.PIXEL_GRABBER_RGB_avalon_mm_slave_read                     (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_read),           //                                                     .read
		.PIXEL_GRABBER_RGB_avalon_mm_slave_readdata                 (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_readdata),       //                                                     .readdata
		.PIXEL_GRABBER_RGB_avalon_mm_slave_writedata                (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_writedata),      //                                                     .writedata
		.PIXEL_GRABBER_RGB_avalon_mm_slave_chipselect               (mm_interconnect_0_pixel_grabber_rgb_avalon_mm_slave_chipselect),     //                                                     .chipselect
		.RGB_TO_HSV_avalon_mm_slave_address                         (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_address),               //                           RGB_TO_HSV_avalon_mm_slave.address
		.RGB_TO_HSV_avalon_mm_slave_write                           (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_write),                 //                                                     .write
		.RGB_TO_HSV_avalon_mm_slave_read                            (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_read),                  //                                                     .read
		.RGB_TO_HSV_avalon_mm_slave_readdata                        (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_readdata),              //                                                     .readdata
		.RGB_TO_HSV_avalon_mm_slave_writedata                       (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_writedata),             //                                                     .writedata
		.RGB_TO_HSV_avalon_mm_slave_chipselect                      (mm_interconnect_0_rgb_to_hsv_avalon_mm_slave_chipselect),            //                                                     .chipselect
		.sw_s1_address                                              (mm_interconnect_0_sw_s1_address),                                    //                                                sw_s1.address
		.sw_s1_readdata                                             (mm_interconnect_0_sw_s1_readdata),                                   //                                                     .readdata
		.sysid_qsys_control_slave_address                           (mm_interconnect_0_sysid_qsys_control_slave_address),                 //                             sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                          (mm_interconnect_0_sysid_qsys_control_slave_readdata),                //                                                     .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_address                       (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address),             //                         TERASIC_AUTO_FOCUS_0_mm_ctrl.address
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_write                         (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write),               //                                                     .write
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_read                          (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read),                //                                                     .read
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata                      (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata),            //                                                     .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata                     (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata),           //                                                     .writedata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect                    (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect),          //                                                     .chipselect
		.timer_s1_address                                           (mm_interconnect_0_timer_s1_address),                                 //                                             timer_s1.address
		.timer_s1_write                                             (mm_interconnect_0_timer_s1_write),                                   //                                                     .write
		.timer_s1_readdata                                          (mm_interconnect_0_timer_s1_readdata),                                //                                                     .readdata
		.timer_s1_writedata                                         (mm_interconnect_0_timer_s1_writedata),                               //                                                     .writedata
		.timer_s1_chipselect                                        (mm_interconnect_0_timer_s1_chipselect),                              //                                                     .chipselect
		.timer_0_s1_address                                         (mm_interconnect_0_timer_0_s1_address),                               //                                           timer_0_s1.address
		.timer_0_s1_write                                           (mm_interconnect_0_timer_0_s1_write),                                 //                                                     .write
		.timer_0_s1_readdata                                        (mm_interconnect_0_timer_0_s1_readdata),                              //                                                     .readdata
		.timer_0_s1_writedata                                       (mm_interconnect_0_timer_0_s1_writedata),                             //                                                     .writedata
		.timer_0_s1_chipselect                                      (mm_interconnect_0_timer_0_s1_chipselect),                            //                                                     .chipselect
		.timer_1_s1_address                                         (mm_interconnect_0_timer_1_s1_address),                               //                                           timer_1_s1.address
		.timer_1_s1_write                                           (mm_interconnect_0_timer_1_s1_write),                                 //                                                     .write
		.timer_1_s1_readdata                                        (mm_interconnect_0_timer_1_s1_readdata),                              //                                                     .readdata
		.timer_1_s1_writedata                                       (mm_interconnect_0_timer_1_s1_writedata),                             //                                                     .writedata
		.timer_1_s1_chipselect                                      (mm_interconnect_0_timer_1_s1_chipselect),                            //                                                     .chipselect
		.uart_0_s1_address                                          (mm_interconnect_0_uart_0_s1_address),                                //                                            uart_0_s1.address
		.uart_0_s1_write                                            (mm_interconnect_0_uart_0_s1_write),                                  //                                                     .write
		.uart_0_s1_read                                             (mm_interconnect_0_uart_0_s1_read),                                   //                                                     .read
		.uart_0_s1_readdata                                         (mm_interconnect_0_uart_0_s1_readdata),                               //                                                     .readdata
		.uart_0_s1_writedata                                        (mm_interconnect_0_uart_0_s1_writedata),                              //                                                     .writedata
		.uart_0_s1_begintransfer                                    (mm_interconnect_0_uart_0_s1_begintransfer),                          //                                                     .begintransfer
		.uart_0_s1_chipselect                                       (mm_interconnect_0_uart_0_s1_chipselect)                              //                                                     .chipselect
	);

	Qsys_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c2_clk                                 (altpll_0_c2_clk),                          //                               altpll_0_c2.clk
		.alt_vip_vfb_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),       // alt_vip_vfb_0_reset_reset_bridge_in_reset.reset
		.alt_vip_vfb_0_read_master_address               (alt_vip_vfb_0_read_master_address),        //                 alt_vip_vfb_0_read_master.address
		.alt_vip_vfb_0_read_master_waitrequest           (alt_vip_vfb_0_read_master_waitrequest),    //                                          .waitrequest
		.alt_vip_vfb_0_read_master_burstcount            (alt_vip_vfb_0_read_master_burstcount),     //                                          .burstcount
		.alt_vip_vfb_0_read_master_read                  (alt_vip_vfb_0_read_master_read),           //                                          .read
		.alt_vip_vfb_0_read_master_readdata              (alt_vip_vfb_0_read_master_readdata),       //                                          .readdata
		.alt_vip_vfb_0_read_master_readdatavalid         (alt_vip_vfb_0_read_master_readdatavalid),  //                                          .readdatavalid
		.alt_vip_vfb_0_write_master_address              (alt_vip_vfb_0_write_master_address),       //                alt_vip_vfb_0_write_master.address
		.alt_vip_vfb_0_write_master_waitrequest          (alt_vip_vfb_0_write_master_waitrequest),   //                                          .waitrequest
		.alt_vip_vfb_0_write_master_burstcount           (alt_vip_vfb_0_write_master_burstcount),    //                                          .burstcount
		.alt_vip_vfb_0_write_master_write                (alt_vip_vfb_0_write_master_write),         //                                          .write
		.alt_vip_vfb_0_write_master_writedata            (alt_vip_vfb_0_write_master_writedata),     //                                          .writedata
		.sdram_s1_address                                (mm_interconnect_1_sdram_s1_address),       //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_1_sdram_s1_write),         //                                          .write
		.sdram_s1_read                                   (mm_interconnect_1_sdram_s1_read),          //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_1_sdram_s1_readdata),      //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_1_sdram_s1_writedata),     //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_1_sdram_s1_byteenable),    //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_1_sdram_s1_readdatavalid), //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_1_sdram_s1_waitrequest),   //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_1_sdram_s1_chipselect)     //                                          .chipselect
	);

	Qsys_irq_mapper irq_mapper (
		.clk           (altpll_2_c0_clk),                    //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_2_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_2_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_2_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_2_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	Qsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (altpll_1_c0_clk),                                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                        // in_rst_0.reset
		.in_0_data           (obstacle_dist_0_avalon_streaming_source_data),          //     in_0.data
		.in_0_valid          (obstacle_dist_0_avalon_streaming_source_valid),         //         .valid
		.in_0_ready          (obstacle_dist_0_avalon_streaming_source_ready),         //         .ready
		.in_0_startofpacket  (obstacle_dist_0_avalon_streaming_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (obstacle_dist_0_avalon_streaming_source_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),                          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                 //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),                   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)                          //         .empty
	);

	Qsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (altpll_0_c2_clk),                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (terasic_auto_focus_0_dout_data),            //     in_0.data
		.in_0_valid          (terasic_auto_focus_0_dout_valid),           //         .valid
		.in_0_ready          (terasic_auto_focus_0_dout_ready),           //         .ready
		.in_0_startofpacket  (terasic_auto_focus_0_dout_startofpacket),   //         .startofpacket
		.in_0_endofpacket    (terasic_auto_focus_0_dout_endofpacket),     //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	Qsys_avalon_st_adapter_002 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter_002 (
		.in_clk_0_clk        (altpll_1_c0_clk),                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (dc_fifo_0_out_data),                        //     in_0.data
		.in_0_valid          (dc_fifo_0_out_valid),                       //         .valid
		.in_0_ready          (dc_fifo_0_out_ready),                       //         .ready
		.in_0_startofpacket  (dc_fifo_0_out_startofpacket),               //         .startofpacket
		.in_0_endofpacket    (dc_fifo_0_out_endofpacket),                 //         .endofpacket
		.in_0_empty          (dc_fifo_0_out_empty),                       //         .empty
		.out_0_data          (avalon_st_adapter_002_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_002_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_002_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_002_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_002_out_0_endofpacket)    //         .endofpacket
	);

	Qsys_avalon_st_adapter_003 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter_003 (
		.in_clk_0_clk        (altpll_0_c2_clk),                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (dc_fifo_1_out_data),                        //     in_0.data
		.in_0_valid          (dc_fifo_1_out_valid),                       //         .valid
		.in_0_ready          (dc_fifo_1_out_ready),                       //         .ready
		.in_0_startofpacket  (dc_fifo_1_out_startofpacket),               //         .startofpacket
		.in_0_endofpacket    (dc_fifo_1_out_endofpacket),                 //         .endofpacket
		.in_0_empty          (dc_fifo_1_out_empty),                       //         .empty
		.out_0_data          (avalon_st_adapter_003_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_003_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_003_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_003_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_003_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_003_out_0_empty)          //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_1_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c2_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (altpll_2_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_2_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
