��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P3K��$�?~������\͡��dk�⍥xm3T��8�׬����:@Ӻ�n~��6�*ݚ������a4�**�1'wO���?�N38W�'�T�u\�V$_c�osQ��o��5�x�-����7c�­R|L1�ni ���_��Ι͑��Sy��d���c�bm�@n5�~�Q�q�Aź��lE�:��xm�~)$t<~}!C�M�m�3�Kہ�eC����I��aj��c*^L�U����ܖ��<˶�]��9+�������|�M�vy���ݭ\���!�v%ט�*ƞ��❡��qQR?��b��=�y&����_0{�T��CjN��� ��K�c �md������MZ����V
h�v����*��� ��o�|��?Lx��,�?>���d4�4rb40}\D��uW8ʿ�S�\����K���2�Z:�*����Qe\v�PG,��[l�&:��D��·���p�����LVI�� 9�EuS(�'�,w�Kg���![��F߲��1U��a;#��RKYV�zx)�E��4�L�݌���ч��<���J'�6�*k��-X�&���h_�O��ߺ{����R������<���`�K,�� aq�������s��Y�%wy�6֚�MJr�n��6�1�h�C����+�`�V�L��k��̔���P�ta�c]�ߙ��T?N�:+xL�]��tY[m�}�H�N�M���p��k�8v��#=���3Jg��ʈ&��qO�;��
&]S�,�Y��Ϙ_F��])����%mٚ���lF��վ�]�f�E
S1Q�fp;2[Z]��$}�#J���w@�ʻ��'�~�"���K�=��y:�5�����6!8Vّ���XZ3Qz�� ��N��3�G@�!	f]a�-�{ۦkk��U��#D'g1Fjr~�4��lOz,ʞz��H�Ά!�Ȼ�� ����cJ�1��J�\���I��I�1'�#�S���P�6��V!G��i��hO�i��CҖ$�������VQ�\��̔x�����/�W��|ihi6Pmj��u��ԕ��&�Lp[��sP;.���{V�uX��Uh�Z���Ek~��9��=����V˹��
|�]{��Ϣ��tY�������Ͱ�f� U����N���:�������#c�r�\-�l��G�jq#Q*���ϡԨz��~�>[O��]�Z7���,�[#���+���$�.�pN�)I�I�k�0T<�Q�����SәȘuC6(z\�c�?E4����r�mD��%ME���P��1��x�?�d�y����s�-AC�L����dU�4�v2�:�����[\0�&�$�<|������$��ot~gj7q�-M���Uy4v����|ɡȾ�މ>�K�a?�Sbx&�s^��Y�u?	��s}����,�zo��o�jK�y�R�7�!�hy�>vd%Q�/�e@���T�Λ�rw0�K����N?\�M(/#R9��3�"F�����'C�{ ����(X��n�|����c�U� ���BF��87��m�MA�հ�R:���5MD�L�������/��rJ�Dq��СQa@��تAu_2rybx�)���
�rGs$vOn�:W೺�<�2��H�����c���s�'J�<�DA�M��}�8�ٶ]���;͕����H� �g=@��e����"2F�#��@���<.i=�C���J⊯O)!�}~����1�G�x�����gw�b^�J���J�����m�U��"�~�>'.��ν���0���s=����t��kZl����f�_��dB�+�
q��ͮ�}L�ŗ]��ڕX�@�G��z�����{N�_Iٛ���� D�*���fo��͹����*���\K*m��kƟʚ�.��"���j�	����g�H����2���	�A�¸	��̇L`=�+e���+n!����}�Y��O��]�O=˯�~���H�Pݢ��T��'���S&������G�F|�vlR�Ft���Ur��è���^˰�FȺ0��eas������m�o�zUZ��ću��v��~���.��+�sp� ON����Ҕ~a�{��up��"�R�B��Ip2��$�g��L�Ԕ���I��Uhh3v;W���laq�7��!�|�L�=m\������!.ܼd�<���~u���ܓ�3�2�Xҁ��H7��eN&j���&GB
�C���~),tގR]���^,�*��
$b>�u��~!�=T�v
�#q ��� ,��������uP;�[�)���ę�\�����v�{�I�M��ې&*b��v6�u&f�\�����-��*�QaU�����~;Vq[涞�'K_�xt�Y�$�Nn'Gave��O�����4���L��1�3�l���A����|R�C͘/{� Q���Y��+7�3�.�m5��w�R{��DҌ�E�n\�<b �&�W��v7�NɆ��3�?����m��/O�4�>&O� u�f�F�hZ����`�W��Ǟ�	p���O%�<�T�t&R%���#�-��^zώMO�#�gAH&�uw��Q�s�i��U���,y\;_�nw�?�$6?��~����Ü��biw5��:ђI{����O����z��F� ��f�9�+N�(����[� 1%���~�?�Z��_�NR�Ɵ�b���ߥ�L�0(�xK m�X4r�D8s#'�͸�8�������(�p��l��.
y�i_��:���Dg(��D�w��M
�� y���>��҈`�1 ���BS��2g��i�L���� ���k��v.�5�l[D)�0;��M��8K�Ǥ�ɭ��RX��]��#|��n3�J��ކN�����Uk�c�(��Z������T�l�N�3Q�����f	�_����X�2D_�u��4q�y��s������*[�I��Q4j�T��E�<'�bI3�#C~Q���_��&���7���$��
x��G)��- �eHCbDDTX���b�2�!mlHc(ļ������~�쁚�Z�!Y�ɡn�:�5������w��u(�H1��|>��2|�,����^�H�ހ���DwWĠ��D�5yLg8V܅���צ�`٦s|µV�:����z�R�X�������VJ��,3@_auǿ�f�%W��u��u4JnYo�4u��Q����.���>�������ݐu�!���\�2�Yi��n3�.��!<Q/]�"��g���e�����߸֑Sfg��&��` |��6��,��xzjK~rN��b�VCC����	�� ?Ox��u���mg��'CN�.v�\ >�=�gC����E�/b�e��p���
��bœG��5�L*&���6�1����t�@]`����M�se���9� )�˃jHO�E.��`|`�������W[w�1f����j�����V���$_2+�<1��^���U��@¯VAH��+�����Ȼ�!��������ó: ��b_�y�D����Z:r|U�B	,�L���@z�c����ۤ��VK��X�>�I����L�v��gq�,�	&X'2�9��@�h9�+(dM*�&�t:lb7P��fI��U�ʖ���S��rZ�ՑG���E�w���Ձ�D�E�T@S�pb��T-�u��Τ�K���!�d&�<p��+�F��Г����m2��t3��S��8�6ʨ�Lf���)H��q�f"�b�@��ȣ�ϙ%�'�SU�$s�xg_}}v.7�I_�A֋x*��u��%9���ޚ:+�4�� oŮ�K�� nI4EV�y���������x���.p�:�j�F\�C\8a�F���t�Bi��B+"2W���xEs-�`�V�m+d���|J%���L����ڬ��-�"�3�-��-gVi�wɛ���i�/*�og�J��	p��Y��� IuAs�&$�LK6�Ĳ{sҒ��,�ɯ�|�8�)� �kbH�<�N��U�Vk�x�����;I#R�J���'�F��L�0Q�\lu:6 �p)�̗�%��i��&k�#:#����8��y���>�J�l���~[�p(�,	�	��露�`.��4+��r�._Ɏ�5�t	ajy¿7�_���u���<X� �����o�`$���}�b�O�dˠ���_~&ꃃ3����Ǐ��ҶS��$�~���-X�U�e�,���+��F�I���5�"{(�9G4�ܶl���T��yֹYu�Sr�+��-�s(�r�҈�q»,*��Q9�|�������9��
(�q�*Ơ�܊���ō�:G�(nsQ�:���LUl��T Vzx��C�N5��A����g��p��?�1�+6�D�)G4A�q�V��6�g=�o��$UB�+��L����~K��������,���E��4�0���c��!�G){����aO������[鎜lLb+������ӈ�(�7��]�~4��3�B$>�Hb>J�(Gvq�˾&H1V�	�����(�'H��)'��)��8�T5�y�Pr?�O��X1Ǎ���s��1ח	 �@'���[gaw�1Hn��֐��ң��l�`˫���K=dq�b|�G���;��*-�f� �|��Ǜ�o�'��a����;��9����}!�Ed#�͊���)�r襰 ���(�7�Z�FZU�r�: M+�X��X-ѯ�D��JЯ2�!���a`��D���g!��X/�fo��%O$!�ߔ~��*�㔠τ" wD���k�v)(�����󫁰Ǜ 3� qg�
�^���ִ�����#Y=����f����fMV���G�:,	��g���iC��W�%j@4��w��Q�ّ6!��ΓnȮ����P�l�N��ٗωK.��1N��}�X�	�(U�V�y��{����`�8L�L��d�KM�nD}����RT�ښ	
����%�L�E/�?�m%5�A�E� z���w��X��=���c;-U2�cP���/)g3�����1�e�Ɓ��p[�m��Ԅ)&��3���?a�cB%��/��ډU3K]M���Zg��-g�=�,[�nM�k��]*nJ�>Z`n˃7G����F����"+`�)��z�r=d5���'�Џ�Ku0n]�'�O������,��J{T�>���L��/ML��D\�4��k̚���Uy���Y��'k�x�T$'�c�e/��C�%���
O���X�ɡM��d6
20F��5K����
�1x;����{9 u�i�䅪n���::�mK��W��Yh��D5����VK��h��O�M,:�\�m�69NE}�B7z������q�j~�
c3�����?�-��2B�UU���zT��F�4���n6��D*�(q$k1z9�:7S���qW����L�z)@�/���j�׹T�(�^'�Eux�8���:��2q�D���?�V;�����÷�"���i��G�AR��q��vB}O�D~,{k�d��ǫ�Qrl�<UE���}q�����mVz�~�,��Ҵ|;�8��I��Ǿ�\����B���y��<����}�4M�!�g�z~sF�G�YC
&��v��m���BN���t��bj�֚6�5�y�.����'�Q�Lv��'D��hZ�Dy����S��Q���iN��Z��ɚ�p�7V��1���dm�&)��Z���	Z��QlN^u�
=��+��_��߮:AK��Ƥ�!�D��zJ%H=N��)6��>雦<�<t�N�1���]��C3G�T�i
��`��N 3��%��vGu�d�����:306pЅ��i�O��5~��گ�eHJ�fy���ΐ�7���H��t��3刑�M�u�H�C ����,��O��C�f�֤�c� J����S��������Qk3˵�O���,�Ț3��S���S$���M�$p;�ll�0�^����F��Z~̗aC+�x��
j�i@��v���L>�&6nBYF�Eӄq�`	�ގŃp��5���j�q�;p d��.�9�w.n\��5훥��"�6>ƙ�7�*����H�N�Ȗ���
4_�^ a�uf�S;���$c�L�$�+u5���'�It��\ͪC/��%(�m:�NaֺGkE��A��Ar�<���]"҄�f䛃��[��O�2N[�ꃤS�X��%1$)�Q��V�E��tv�Z�| �[�X��3hq;�������v��� -'_I�_W ������+�m�"ɟ��T�+��I��}D}r�-��:�o�긂_ͳw/�K�S�3��Ɇ�<�/���
%���C������4�H7����y3��n C0���T��۶�
W�[|��;�b���� ��9}xDl���{]M���@��a���tx��4%�Z�D�� �b���!MY��L�_��6�t�;�ٟ�޶=U�7�Fm�6)9k>b���Yt�������tKwl�Yָ���Y� ����#�Ȯ��3�~ޅ��Y`H8�J Ɵ���'+`��r�g�o`a!=���$}��\�S��f�J��]b�-��&��}�n�c��b���>2u� "`�w�N�gh_^�	�5�mW��-�<�l�����D1��K>s�!�_�J��U%	��z�W���p~�˗Q�J������UL 4x*�,��b=����]�Jb�7&t�Q��~�������78Y�6G��Ӗ��߈���̈́�G3���	���Y���.E�DLp�y��Z�֜��˦�i��y�5�j������~.����/���@��b�j�O��E)T��h��n�Q�r�)r_nFF�s�Q#����eH�.�1Кs�cFޖx�c�,�U��� F̃�~V�v�������c�#�VT�����iA�t��9��>&��RE�pBa��@��l��6��o�o�J��e3kUh簮��b��%����ZR��v�w��{b�7_xRp�/���;���]��.��^�LJt���Rl~�0M��-#�lQK���&N�ݐ
��a�"��%�L	P��X���ċ`�13�����t���@X�aa�S�s���G=��e�~�u���=�k��)��U/߸��c��c_�b��s�Qc�6{�U�I��V놼�3�f�a�qK������Y�B�.�gC�m��m�/k��/�ɛ�8$��j�J���;�������'k�~?�67c��
Vtd�_���n��]��Ӈ�9�|�8�5D�+.�W
Z��v��s ��w�� �&���<ٹ:7��O��[���*3�g�CN�-��z�*O����Z�� �K���l���������]���Tk����}@��=�S�Χ�?)���p�c�,	Ѫ�|�tm�ZwHǥ����b�.Y��=�o��إ� c�1����.5�L3]#!Nس
x�zd���u�_1��6�f/_���Lj�2���-�Ȭ>@�x�/���Ú�r�g�����[G�h�g�x)�O�ư��p
�;w ��/{	��_|~�~/�P��]}�([N9��`�0-u�� G#�## U��CD���G���^-:S�Km��S�n�{Q?)�N��U�|��\姻n�ʢ�BV�����+��Tdo��Ґ�5��r՚�ۮ����K���V�Ң�^%C�dYT{SO�xIvX�d&��ڨ:�ypn�]��ܞ٩�/�H��tJV��;:ËiU��d�uPe���7ɉ�DP�~�1�V��L{:�Nju���o�0q���%Ѡ��`���|?&+��n'�t|�Az�z�i��@4�L�m�>����:5Os���<�h�3�~�!Ȇ�[+���n`I`��?��i"�Rr��:�-9l|���P�ƌS����r��X�;/'q ��33���?Z�L<�Z�w������1��6K�#k8I`��rp϶7D�q��cK�uj���E�G&����&�A�>��Z�J�pz�����
I���2���X�ЀpO�r���ݽpE�;��H�[�g�5ٞ˟%Y�l������б�R�j�
՞ede��1`�!2�Evۈ��*_��' ��4;��]�C~��ڐuw���y"�rጫI�	�W.�;�X3��+�C�t~��[N����ؑqÖ��{8�6��A���b��}�A�z�(�/ɪ:j_�9���x�l%ݮ Fsr���}������
'������İ�ÅUJ@zj��r�h����L�R���9���r?�;���s��,���ņn�$��J�K�\|�]�>0�HCSkǲL�r�8
Z��&���{x��4��R9�$���8�Y���.d�#wJ�)�0����jm'KhysM�Rc�Z��[$�+�����&#�~���6���$�QZ���p�E�=�o5�)�k�4�`�L՞)�)T�Q�a���wb���$�QW��Awb��sR� ss���v�h��m���+ܖ<��29�Ы?��P��շ.����Q��}�q�z1�&��8cR���7����{�>>��Q^V�4yG#�V+ �$��}��=��Iŧ\��6�e�D�`�/w�U��Ъ7K$B�
1�;�&��k�m�D��=���5���g���c޺̜Q������F=#Nh�:��O��lN�_6h�X���>��7	+�=����m�HLP\�"���h��}�:��W��vk&0�xpJ-�Խ���e}yY��7�B� ��(��F~\J������x�\�2gL�U�Bx�$F7��t�E�$M�VA ���wa�ab ;dr�\���W�RK�8rbk֩�%��xgDE�T��3R��D��l�}g���ԯH��is��Z�Ճ3���Ȭ;�&!�:2�#L'-� ������~yO�l;xP����@�l��0E��t���O��V��G�U��2��+���9�ދ��#3�#�R�A'�F�ڱ�'��z 	`����A�g޺���"�]#1=�Z��vP��?Vz20B.���	��PʫUD���~"7�q2䚀ɝLd`z»r/��{�e6��V�YF�6:.��&o3/��#QF��[Zg�+�ޑ����(Ȼ�Zf,\FE�%��~q���dĻ�sx�餾��H���V p�J��W�� ���� '�aB��#�+49�_�"�f�@�-����ofj{�`��Exa�X���;g�Ɩ's�ݗ�q�v�Oty��-ߝ�JU��K�nZc��e�:v�ۢY�&�xQ��Ȍ^�P�oը$��#�Db����󉚥��4�6 �^�s��sѮ��;���_���R1��$��E{�̧?9�fM�֔Nd��3-�J�%@'Q�h.��[���,��GGk�P�t���0[x�'ǣ.����`<� rF��-��lw��d�*.U^����]G��2�*��U������^���y�zA3lrZcI:�,�O9�W���E���`���_h04���(�,� ��5*߹4�;SC�m����0�Q#������t��x(��p51�p@����*�=-�A]��&���e�nu�|������T,Q"ʆ��k��S��k{��4�߶���̠�BD� �
ed[���QG&�Ȥzڢ�.3h���r�T��R���[hW��1�я�tn�K§>��R׋p�S@z�j��ty]"z�gɶ�,�m��
I�#
a+��1��Z�Έ���� �)�jg�d�qus��7�syQ�YP�(����o���׊�ZX��͝s�|F()^qJ6M(��q�X��d�*N���j���6�o�j�q0\�J�\�����7���P�ݨ�P�7�k=��`��Dz�롲�k0�Vm
�������G���[>�t�>2�Ǖ�ْ�U!?O��}1�����vP{9>��,*�V�Xp{���a�N@��v�r��#?쉫�,�Y��a��b#s�}���,�܂�"n��w>�P��ʺ��gʑ�(��p�F
�St�*�*l#w�6��rђ����H���F������|6q
�08�A��A_�p��U�c���_�(Y�5�UV,�T��P��S!��U������d��j���z�/�.bY�?7�}�BSu��Ц�D������N��%��@�m�X��"��	ےR|��b��B��xyo�r~���N��?*U���BÎ0�_��pps�`sV�%���l����7W�*�S������[����
�X��`�; Ɗ;F��Z����-V]���4;��߂�~�L]m@��y�:�I>Wae�^��>����.�tNɔ���&�-��r��[O��<���#��f�+d_��NR��%WR'B����$��sd�y2Ņ�ԩ��N�����sv6�dQ�U�Lsz��=�%"�u8(�+���u��>�]4�FM��ä�c#~@�6��X^�%9�o�%:h������[� �@���[?L�|�M	T��SJ磢	2��\�{�IT�_�;̣X���� pzj"8�p��� ���d�µ{�,ӥ�\?��Z̏�9(��Ј� w�i+�T+��V�q�=
�������yCn�JW'�t�Ӣ4R0{���t�����Y+(���f�r&�s���Q��)PȦ2H�ə�blu?-\Ε���2�H�=J\(|)������Gx�^��e;����ö��e@l��X�YV��r�ʽd��)�ى�74����5H��� b��rY@?�BY�N��w��yGc�N���MR⻺�r�ʡd����}е�]E%=n��y���-y-L[i��u���w�� ��fa:�|b��U$�";�y����B�!���R?�|�{��1,b/+�=�h�]"i�`��`aT,�bɖ�%�K�Nt������$��صP [���\}�y�݇8��L��=
�<

킄�>��Vp�mC]���=/g���9Sm�L�(��h�Y��HSl�"7L9���듰�G��d>�5a������@��z�>��mE��q���!� o��B��"(�y<�%%�r�ċ:ξx�q�$E|C�V���M�rߏ3=z�iQ���<��E
� 6�H�JGz`��3F���yVղ��VU�B��� �@�O�U��^O傲Mwv��/��k�����y7U�HjA)I�v�2�'*f����T��[��|�gf-�Y��ߙ}�4�B|q�GU�q�~��6���L���&��NܿZ��1�M��N(uXS�/��h��x�<�ɀ�mbol�Db�%B�x��_�>�{��K2��s�f#�C}���rު�0�'��ޖ���i��>�}ˍ�� �+}g�}׮�W�1�{ò�2=E�!졓F���og�1��]��M_
�Z�PK(��T9ȫa+r@���T{b�3��	��EI�O񢰪c����pb��I�=�&�<i�+4\���D8���4:�78�U�/��K�x�o����Ji�VLS��	Qw�����A����il&��pa�V���k�5���'��`�0c���T��Z��Яrw��LO�]] �W#�3��r�WyM�[6����Y�`��I�/6(����5k����R�4����4p�W��J���rw���%�Nhؽ`�E��qԡ�y����w�F!J4�C�.{�k���_���%���s,l�ǻ��run�
��x7Em\Epjw�\��Б�8V���^����Gꆤ�͌�ǯ��n�K,�2X�\�<?;1���k:�5k"��Z'0ҥ��x�K~�s�<o
֎$�T�����H�l�1U��8+:�^(�K7W��JC'����?��O
���g�M�`���T<��)�+-bmB�l%d���L��ظ�U����!�/�O�D�ݾ���B��e��r�M�O;:x!jS�DW���d��.0�V�]������+�K8x���\ƻ�o���p�j"^��T�y���_�I�L�+�!��20F��#~�������k�8�$��j|k>K�����W�XC�?eL��J,F�k��;<�':$�����R�N����������>���z���z�K�kv�{��4�l�sN�
�ügm�<n��o'���? ��I`��M��)1�# C�Ky-�Ӏ�}�6�Q�P=�  Ѳtp^��r�GPRfGջM+K�R��_����q���y����4|	|Ej@��r;��3A�sZ��XK����~�'��7�9���@��uR�P�)��������tc%�I�K�Ȇy���D=�nq~��iI/����,bt�"��/A9��{�z�\���������|�oU5��r.ƣ���aw�PZ�4U}�&�Z�*1v��dݩ#E�h�����o�0t��h��̢����R[x�e6��&0tZ�s��ӝ�`��� P!1���Uf���`J?'	k�6teE%�bA�9����)�j<4b5���6��Z�F�y�NVM�G.�����ď	4QF�mS.B\]�����kPN�0bq%�0�}x�vɃ=�6�*�єd��Җ�]q��k�k$��v�w��`��Ǯ���z+�K�����۽3ޑ���-��$E� ƹ���8�R�Tb�mzs���]�W�V�06}K`~�D��_�w�wǒ�̈́��KzCǊ�����52�]�o���/)�bjh��XI���}�U`kӜ��+��@��<�U��.�a���+�����4�aq�să�X����w#rih\�J�C#����z+6f��Dg�ۗ��Ë9�p;��@ ޞ{�Yy�7��}����so��vg��gb�0O���*Ț�w�l�(�㶊	���ћu��*�����w�F��շ���zs����H�K;z�����g��:��uJ6���0⻃�!��Y?���{?�4�F?�1�	*��\`)�(�lH����5*(>�����K��ՔW�3��8��*�K��}m���m����s��1E��j}Ib8��F0ycQ�R�ͩ��Z�b�;�kv�zW=��8�+(�-BJc��甃Q�	��J���ds�H�n�1Y��"l|� �o���'�tNX�4:�MC���2����y�ח��r����Ȟ��@���H�m����I7G5��Z��k$5#k?�����i�@��x�͑��l>C���<����U��+
țc��`N���c�����ʤ ��>,�ʩ	��:q��x⨭yYa�boYĻ4��L2����Yaܪ�>��Sڄ �o��M�S	e�����:b*�!
�|����"O�����P}$�RK��]u�"��?jи������T$��.23���R����B�@���Bv ����/���9�mբ��bU8���M]R��c�L(=:����yXz�����z�h��7b��à����/���c�ɤ��K��fRWЕ�BXR��	�ި5�89"*x�X��>�ƔY�i�6�G��7�bL/�p#����T]^ѵφ��q4�4�T���*��J�r��
tW2"����'����b5	�[���ʛ�ѡ�	�
���~�o���н���w^�"�Uz���y14@�P�G�g�5��-	9�?8׈��wV��~�&��~�p��o�1�M[GpX)�hL`PF�U�%���|(L7��L�e���~�Ǜ?âlo�Lڲ�!�Ϫq| �e��=���$�;; �P��9o�#N��ZW���Ă9�n�v���o/<YU�5sm-jun+��O�]$�\Vy4C�rR��iH�c���H���w������`-�����O&*"%t��Eɽ��Ƚ;������+�t*L��j�`�|:�_s#�ڎrN���y���M��s�=
��NV4vf�_��@�5E[��L�.x}�L�C¹��2go�1,�����)Z
��̰�&�R��\��X�-���]��rl
t�؅�����Oy�^��24��*�������שL���ڂ9cU(�n�-�<�����W��!$�C]QLyDC� �C:�Ӛ��s���ğ��.����<��0�E���$�,� �X�ߙ���Sԑ�q�UCfF��urK��S�urÒQ�/E�Br�s'?+N<�	���UMe?VR���gH1<��Z�` ��f[}���:�؁�KL��,@�t�Y��Q���hlm��K����ն�����;�?�1���q�9���*#�]�nKge�ϒ�a_�D��zp�B�`��S�|;����Y�LەS�-����n|}���&|�RP�+u�Y��u�=T��²���?"Gw�$ �Xg���p0Ch;ROy����6ޙ�ő~}^���n[:Rk���