��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P3K��$�?~������\͡��dk�⍥xm3T��8�׬����:@Ӻ�n~��6�*ݚ������a4�**�1'wO���?�N38W�'�T�u/���~Wpm�ك>K��]�q�HI��w@��t�hB���"#s`��	���c�"�9��X9��(��ʌ��lr^��V�6�n�!Y%����mkqA����Q�T	�r_�Pr���������;�D�(74J���Q���7=~_����D�?&�����J(L�ӯkc��r�Ɯ
�MR��۸H>�Q��j�7>�/LDӊe�	4�ѳ�ʗJ�/|?߳�J� 6�L��)��kgá��'��Ȕr�R��r��n��n�P�L^9����\�	[�./[_�텗n��u��!6�U�b�b��?6�$�
��1.t�h5z�3��4�+�B��b�@Z TU�e�8����kWgP����I]qvA�ȸK9��},��I��L�~���ο�x`l�4��gB̪��n1 �.�}Fe�h����0z��㤳�s����,?��I�tk�A;�0�9��7��ӵ��z���x�3�\d���?vcWkf�F8D������8.�����6���Q�l���]~+;
~�J�⺑ab�?�q� ��+$eH�4T�+'G�F�i �(�;.
��'�	��'X��TE��B��"�ܿ���.�)�]`�Rv?�(]G�Y�C��F��C߬b�=1#�u^�EB��8_-��nQ���M3�	>q Sp�3x��yf����O��8狗3�K�+&\�_�$b�>}���h/�����z�s��1oKI���W������N����$���3�J��O��#����&#��X�keF��;1-�!�����&��'� OK!�Hy�=�]E=���(c���	�q��[�ϓ��M�_��5�]
�_���@�=����V�	j�j�Y��8C����Y��Z���^6�%u�_+N������7�f"]�~�*�@X��t��1�\ ���D����"U��L<��$��B%�?���`v	2_C�����%$XV��aK��5��s�� *l��5&����l�F~�}�����X��jJoT�P@[1LG�ڒl�k7�g�J*���/���WqÒ-,R�]m6�}���V9���P��1d${�o�\b��Ҭ5$����4��cF�꼻�V%�!Ѻ���s@�)�{i�>1.?dE�$=��^^�R,V�M[�r����&&�����Fz��V�4�C��Ʋ�\�N�<FT42$�]Y�֊Gl_XX[��C�ģW���C��c�X���&2�PI?���D����ShIxEI���v/���p�]��B|[�R�6�D�ݡ�+T7Fܷ���yP?�;'�����?�Z-o'כ,���'nե�4��^%�a�Q/i��@Wu|���؋"#	�e��>�����l�aN�����\��u��&i��5���Vo���Y�cD�LYL2����UN8�l����$&����fH�Pib�hyU�x�������N���S�m����Ѐ�9�7KL(ly�,��g
�I�{\~\b���ޱA�H�����Wـ#�WU�uY���y��F��QF�_	%�D��!.��f�{L�I� k�l���[Br�#�jnۍ�=��}���;Eڰ����;{��V���4���x���LOMOB�UW�/G�����L�m��b���d�.+(�[�ߙX�ą-��Fry�MO�}�;G;�eUo�	������b>�>@(4؇Ϯ���X�Vxl!��J4�W��:�F�\����ۈ�>~w���,�Gd�|�"ӷ�˅x��"!��Y�CӶ�_��!d.~���@�n)��}�=G=J�Jg�A�Z��Cŏd&uC'g��vl��zլ��i�fq3b��=�g��\�ܛ���cA��,�{�\ґ&)��=�zxڪɅ�)t�Ǡ��� �%���َ+=r����{���x�~����Mk�.�*����;}�T/����RmIp ֥��J�T�|x�l�A�Q].T2�Lq炦�y�h��qT�V�[��x�L��缹W5��Dԗnb%�6�Dj6�J�@C!5y�մzC�����>	�L*|fR9�G��ϬL�p� ]��OX�
'tP�~�I����DT�	]Y�hD�m[:�5����.����s��Kׯ�I@�R�V�,���A�j���S��s�k&�+��pӗ��MH8�'|J��W��2
=���.�$&dCA���� rǣ�I�L�R7C���r�`�凃���U@:���Ri��>.�{^"�W	�牌������`�9Sm
�����r���U/BV
����&�d�Π��s���
�[8�e�A"�\��]˟^����_�I��K�8���erXI�
���{��4%���0��n�d�E�L� ��� m�t�吴�GM�$KxP��t�y$��o���&�Y1�4-��,ȑ;��h<[��k����1�U�F\|��/32.��}���ny��h����A-�`L�s|u-������9%ǟ(�H�~i!�a�y+Q�"�b,��esk�E��o����j��/�ӈM��S���YN2��:I�5��Y�4D7}@0ȉݛ�xZ;�K��@"��5q��' /�&�D�:$~�Rz)#���
��h������f�Su��3�܍RST�gͥ��:o���?򡿐��+CG�B Y吁w0=l��
%۾��:9y�����ĺ��K��9���Lz?��i^$w��L����<�(<�,f#��;:}���Ӳ3��nf)4'G YDN�B�E8��'��w� ��F���
���'<����T�%%��	y�7�[�芡(U��u��O�c�t�Z;�HGL�^8�21>�����.��3P�N�OV�z�֔dg�g��uP"�=�*��U r���Q3�irۮ����d�;8��� ��7���P�����w���F)����,���{������H�h��%��-6;h"g�p�-�@��Mr�X$�;�\�s�4$��oCR��U�H ���t`4��h�`W3/���j攣y�������8s"g�ю��ҍ�q�H��H�U�R�˃��`TrȄ]������C�k�0��ϧӾ%�=�?��!���m�t*(W�ێ�"��ڞ�]��e�i5Y(9h���w	*Bg UA�2�Ƒ5n���`Zn �
��#�����-d�K���ٗ�!ȴ=YBdؗn�?�HiqdT&�GK�����S��\������O��A�HNQq ���0��𧥔9�٫�[�k�P���l�����,�~)?�U�[Jh�>�@-bW�
��x����"���7W��t�e-���rN����8W�ͼ�&����RY<���'|yLDc~����ee/����K��ϥ�(�VM�F�L�ذ@�e�֑�y昦�$��w�m-�H5@#uT�׊�7V�`�wow���h,��ۚ��[t/����ǹ=_�]��1����p?{M�eK���.��G;}���3�=ЎgUD(��)_�[$8��'����׵I�U6 �h��p ��h1������㴻��W!�d�bʍh����>��-�D.�f.$`���}����)�ó#�TY	�r�D�<��1yg��������Ǘ����^ѿ<+�q��܊W�@���������m�~W%
��?Ҧ5O\=c��E��^��d� �ߖ%Ӣ�Ad��zĬ����q��%o˽_G<�� �>�O���e���R~�ȑ3ꖭ���7=3c��q��F�|��pBѐ���aM�(h���}�TK�\��
�Ӳ� ��t+Rc,�B�b�pr� x��z�a.�C��I��ǁ[�^]`�C�AF�0�A�i��0�1b7A__�$�9�6iCcx���-g�ƻ���k���;����$�N�J��0/��������g$���AP_���ĸzQ7�c%8`�Yw[��m�B�����ЁC��yŌ�R�|��%1oȣ�+�T�qD�+L?�<��wa�&�V��h�%��PN��U��AC0p:ɨ�Μ�O*M����l���|��y?S�h���@�E�<1Z$�?��W��~"	ٙQ���.�ep�j��O\Wo�_�i32��"�(�m����;�`�Kise�X�/�u��d��Q^����^f)R�`�:K���B(<Oyx��aO��k=-��"{�ֻb��R|�H��}сr�uv�q��{Է�^�<�ͤ�߈1j�9�S)���3%�-[0S��_���?e]<��I���E�%�ÇLU 3g2���$��?o��X#��k�/��ހ�&cD��g�L6q)"ý5��{{Λ�q�8�
�����Y�18�����ڈ2a"��9����x��XQ/�wJ	��Y*[�a����{Q����۱щc&����7�B�]����Ul��:�R����Ѓ���5�Fw��j�~{��HcAi��G�Ok��C���#��f�W���۠t��,��70�.BE��RT}����=�O���"�4�;��Rf7�{�@�l��ȰsM8�����<�5���1�Kέ�Y#K{�]��Nu�D��7��({냌ưM���a��9�	����O:p�0� |�g1��gZ`��+@�b�?VU��v�@ȁ��R0ˠ��$���k�9u��J͡6{BMҶ����]g˜�#<�X.�p���X2������x3Kca׃7H����� ݎ��@]I���gq&���,��$����cy����XϬ>ղ0���/"F�\Ʃ٦���eFG��A�~�Ws�]�4�52Y&�B���;Ḃ�i��O��g8��<���zP��}���~Nȩ��4��;۵3��C۽���� |1Q®��(��B���u4�*a����.7����%7'��O�e(ADփ>�r�
C�p,v@�F���(�U��"�a
%�?����?�y�a#�*���^޽Ω�=����B��y�E��r~� N�<�n���_v�g�+J��TB����6�!as���i��]�v*�uȋj]/������^u$�ϛ�=��@]�qJ$���j�O1���f�>��B�@y��؉>�k� �Tҏ]���+�w7]>�B�-㷚��p�1���g��ŖK�l&���-M�(`}Sc�`bYٶ��B/7�}FI���a�oN;۩����Ko �TCߦ��&ٔ*�T4c�	g�x�Uύ�� a���Y����lvE��x�Blԙ�f9�XB�В�L�y�i���w12��El�HS�Jx��U�`g( l���d�[���)ش�͕�[_�-�)Lm�%�Z'D���U��M��`t�#۟�2��z�G���(-q�Z?}�}�?��A��N��7I9U;�^�R��q7u�=
�y �1�{Ѥ�CSc׃(��)]��7�h��ދ"�
@V��1�A�S���>�:ʞ���E���y�,��~���]7�>��6i� �L�5y�����& ��5�d��bu�V�0�t�N �[�@���^0A�O {m+z�hw�����=܁�SrW_�4Auƃ��i=j��>�h'ye��3�Z���U"5Tu`�Y��pg��Ifm�� ԮXa��o�N*�dg��+_]����t��C������iϣp����:�qo��M��ɗ3"��1����r_G�x��RJ]hW2I�q<B݊��vcĳ���3�����9d����M	�Jl�'nm8樂Ϥ-���.KI>��Y��17w#��oT+����>��W���F�6��x���J��@�q9MHbB7R�T	�>���Y�#J��ĳ���f�[��6]��՝�a&#�C����|P�x��);p�g%g��cZF�c�$#B�kk�m�|��2���rwv�Y�G��
,��E��%T�;0�2U�2�C�Ƹe����U}�!���M�S<��/p���-��=|1�f9�!w\4�?��Z3$k2Phd�dggY`����7�K<������x�C��.��m/6D\d�Þ.��:2K�� ޱm�z��m�vRB�V@T���]p��ٞ�o���u��.�Y�����:�$q��V95����| Xl4 ����ܷ��V�36D9D��'b�ϕ���@U�.tJ��ֹN�*qL�i�R��'1��Ƣ�Z0��xk7�(�O��ݵXw� �$s��ը�j��/�q�f�#�KWP�����c����D/����{��~��d9��)7	MY6C���[�0����.y$���h,ɎǍxX�LL%��<�J����YUD.fj�uo/�FatA[�>}:��bQ�I�����1뷥eo�KT��n�h�fz"]�0v
��%Pf�s:��Φ�
;q�����zWOV��#wl-���R�\Vc݃�`i��9Q�ZΚ-pl]���R����-����F�m,��L6�ӳ��Q���G�+G>��m�����Ȣ1�Ҟ'��FǪf׸�LUh߼����������GN�<J�'~��~/�Q�[{]Iv�|ϖ[e�2Z=����#�©-Oo
����^ܨ�gx���jX���6'��}�"Y�*G		�-�A��(!5�%)��Uax������#1�� �%��0o/���ۧ|1���㿰��s�,_×��u�V\z��Z���<!��a��]C#���2��k�����/Rs�P��ᢿ�S`�}�볁��2R�9��H��F�H��g��,�p��q��ɣb�Oi޴Nv�=��`�5����YdSz)?M�	�,����L)���oƐ]TfGH|y��,��ڐov����:�n�m*�[�=s��oUמO�b��Zg�GU �ݬ���'�2���vo#4���-���y�;�܌�q.+�ۭQ|A���у���]i��U��vSE|���=�LHIAƁ,E�N�H��������33�w.3����S2��� �\�W�ɜ������sMi�� 1���Y���S�;���R��E����i8K���fMڎ�Dq/�=�[k�ɕ�X;Z6Z�ʔ���T�"܌�l����(L5�i�����_[��D-� VET1��+�댰��puk'�Һog4�q5`����ֶYA���kUl:O��U����b���e�;eVީN���������9�DKd-����]v�D�êr-��UY�O��W���Jʼ�nH�_B��ހ�^^]��U��x"�߰H�*J��Gv�L��-^�'���"�SA-�Zi�ͪ���x-�\�FN�ϙ$����	�J'��z�<�󾆜D���:�N��)􅏙:Ͼ��X߽P��V�'Zp���<��N��Gu�eոk,���]����/��6�~�ʫ������"�cV����������?r�i%�-��~�[�2��ekq���BKP����{��S�s@��hT��X�"g�t�,�xrI2ÿ��K����9��?�[hLh"����f�ޢ����p"�����ZS�nV(d����H<6\�+)z�ep(�^�P�����}l�b�����ch|X����'��������
z���Z=�Ԁ4�S�?P�VIa,Yڮr��@�8;q��\k��p��:8.%��َk��I3�#Սs1�� D�,�����RD
0���Z@���"'z��YH:�������zG���.@��ngƧ���x���@�b4���ټ��XmW�Ň�k�X=�~��N�O5�����+�e��j�F�Ф��RL�$$�v*�I������YC��x���OW�Ȑ�F>�D�ۿCw�-~Swx��R�)��A˧�H=��Ԯ�7T�>ΚԃS��T �7~�+F��o��5��أ��]�v�3%)�����my{�a$��,~�g�О��vx̕gFrLYz�/n��Ez׉
jM�<v8���퐙�	I���T�H�� ��}83*�Cի<�Jz39�C7$4r���i�giH��?�Xu�����ЁB�,���;�F2�T�m���� ��Jc?W�I��;��=*uW�� �CYS8�{�03��"�h�CNW��V�u����P�q?���4�9
y�a�N���B���7�-�B����.�,�����9� �W.�<1�[E��Li�5�vR�JtV����u��=��m>���2�J����7����!���8Jj�'��XN�H�������t�/���lB�F|�qS:r*�.�L�/�)tU�o�0�V2M����k���V��K�6^>+��w�����yE����8�n��DĊ���^6?S�����a�z(��9L���4Li�Ø�#୻�):%�n���msLi�;gR���Ó�'Y��U�LG��Wc�#��9�I(TC�⡆�db�i>2� �sm�W�R_���"��WG�86�� �������O9�A˚N\���3WJar��"�>+�.��g���Tu��KD0'�a�늕`��C�S�h3+��������*��|g�*�)�����Ώ"��	8q�#���!�S-R&
$Dui(�}�;Y��s/L�3EjΓ����l��#�Ă��b����> c
nLk0bGv�Lc%���`���g��D��"W��kq!�%#�х�օX<ڕA�ȿ�+� �����F0,q*�>�42��]�MZgŁ,,v>��j�2��e����)7O�L�+U�+�Ν1)]S����@xŉ���(��.,(?qq�����n��@F�����E��b7����`�9�Yk�	�p��X���$��e���+@r��3H�>�9�^4�������Gx�:δL��Ǹ~n����d*L��Ua�p;ɔ�\�[�6FF`�P���e���찭�|��zP�A�%˻vZ{j9CD	y�J��>������ f ����#��nгL��S�5���Hڸ�BT��)u�h���J�<�`�f3��0�nA)�绔c�T������ϝA��7�><>!$������+��?�3��@5p+�h�e>����Q�if�v��G�';j�B	��0ljC[#�l^�	T �~$Y?ð&Qp���P�
�-�����[�NM����?����u��������>N��~|��`��i�P�s��&������2AN9z�R�w�!�"I�H	�=[R,���W��R ��}��z�����>�Eo0��
Eqe\��,5�S&�ێ�ˬD��~�j��� j�x���؍�����m
�0���j�N3�&�L�2�h?D\�Gb�	��w����)�3��pD����!�6��?I~���������g������hui�H���<�"�_�
�ǽ�I�=y�T#qg��+�bI߄�7��I6�{O&~�<ڣ"�N?F��^Q���rU��zdhSK�s(>˂��K3���
)沆{_g�3'd{O��pR�g���!�UǏD+��7��M8�|N�i��B�<�_�K]�#��/�g� m��� :�N��m�G�G�����T9�z�V
�t�d�s��S�a
D�  �_���򯫟���A����Q ��`������J{����_$���Ǵ��g'G��x�p����+����It�;j�6{���)�̪���^��q�~���$$�mD�N�1$�J��C�|W�.��>��b�] ݒa]�<��  <�S&�p��h'��\l<�e>�7;|��GMa�::��V��y|�N��d��&�`�"�&��)<ũ��_�ڱ�
��O�Fou���r��7�2����NW_-$	KBJ�׾��c��_�XP�I'~���x�<�1�������9�+�-f���ml����p����(�,f_�C�0TY������.p�t�5��E�y�]��7����й��F�i��w���o������֗;�A�S��2�c�w4հ�|�,��|f|�w]Eo�����=<�s���֕lS���g���{lw��[��[�l�ekr�	��SbX�b���	2qA��01�x7��ʴ��gFM����E��o��h�[K!�|��G��,O:�u�F��!����k#�\B�ɉC`'��f�
g>>��� G�Ya�d1�T�D�d�U(���nN���ƛ4t59ex$n��|��y	��7�C��ݾ�}�~�ֺ8t�*��xb�!�u3F,IQ����q�{�軁?mQWD����kIra;�
��!�)>b�X����� �x����D_���8I���hŝ�s���g�q�-�/��{��CU���Yvp�u=��vs+�m�&$@��k/(���Sy�5���H�� ���p�5�sm�Z;߱ɱd>u��Gr{SС�$�G�<��z�t��������P+˥yi'+���s/I;��tvF.�Q��_Ycqf��}�&�b���s~ �)w��k�0�C���|l�-�R~e�9�~�{�Z
F���V�=��Z�u�$�#4�u��-��7**��'^.�qɎ�G�Ž�
r�tF>ÜAu�)�6ST�&`��A��Y�MʉA�	F��Yo��\p���wCTcNᵗ�=!"7����������]FƓ�{B�@��<�!�m�z���UƟ�.�5�N�W��T�|����X�E��՜� �6�H�e�$��؉���}ג	�� �pF�86�6g!�Asʎ�(�����Z�Fb���;�FxA�3𹀆�. Y���]�:P�
Z�ڗ{%s,���&\��zO��ؠ�n(��5��f�� 1�	}]`c7�Ȱ�����؎�����mce}d����l��ʧ�?mJ�Df���O�!����o��۶�nVA+ߐ�Sp�O�]�N�g��I���e �E�i@�Vx���O°���f�O�Uծ:�a)3� �4!N@/��ͪ%UA���e�A�e�޸�nh�h��J�ww-D �3dT������m ���l��+�~�ߌ��Ԡ,Q$H(`�dJ"��E|�;��,u5��9�QC������/&=�.�z�FvT��S����ls�������qk����|���4b�j�.����͔J�y2I��)�
m�����g�e���K89�R�7����'��,*�]4�WWj�8<�U��Z#�{�&�Eϫ�7�Z�,&_�H'��mk�>mށ4�Ti՘�Ĥa����-�tuo�@������t���X�K�^˔;
HC �1NM�[CT���<{�@�݊/�����]�����k<�
�I�}��؝������$́�𑅴M�b9G$�����0�;5�sou����a�/�P(f�d�3���̀��,K��k��'DW)� Rg\P�N��quTgE��x����f܄<���t{�mF�N���t��>G�7��/m�c;ip�:����l�?��:������1�� >C0O��z�S�9���fn���h�1���;�</8H�G��b�^U�٥w|���]�*ir`�5sp�V������!t�A�*�V8$�c[mA���pmr/�d�e�/�^� �io����Gk�ԓ��K��]`�c��d�V�i��'qtz�>p I
TB�A�o((Y/G!8xX���~�5q�\<���r�CR�}f� �,j{0�~r��ڭ��H���|���'q���d�!>����b�돫l�H��u9�M(~+�4�P	��3�0��i��N�#�������Ց뇖�	rt�ڄD�T�y���3�_u�=>�8Gt�ך�GtlQ<�l��U���=-!M�(2}���
f?���b��,�2}�>o~�{��Rv?�Ә;���P�r'V,���g�CC��hvPzt;�s6��<�.Q�����B��~5E8�B�Ol�(�p��,K�1-⮲3��N���M�OfO�zW��ڨ�*&��s��;�	�Z����c�Uａ����`��fkM�R�u'h�� �ilN����AnVr5��>/r�彛&P��Pq�eS�W9�i&N��a\Б�Kh��c��h�Ai}���/��-@�1e�p��ڸ�sδ�V�� �@T 1R}Ź���E�x��-s��. ��Ӌ���5"�\��¥_,���Z�')c`���
�s����Ka4�����͡"����͠v�օ����=ƾ݉��x%A��lE�dm^3�=t�BP<|c���6=�/���Mo�~Q��1c���x�9ό�H-�Y���EQj�(� �b|��9���!o�iڊ���h�������/筢6K�@�\���P(�,2�fT��V����(i��f4�����T�6̲$���q�����j��û�Z��t��Xֻ���Ř�>��o�\�M:d!���}�k�ڭ�O�߷��v)8�	 $�E��3�T��uuD�����D�Q��]i	�m]\7�e�'�w*W%Se�P�LX1����g5��|��kRZ*,j��ׂ��jA��AM�$'��Խ�}�X�]B��\��[-��hÜԞ*H�W��\/%�'M�<%���n�t�3{Z��%Ux�Ri�4�p�d в�U�Â��kQ{;�`4_U�"���y�	�y��r��:�������_��@�ƈ�`��3~-�[��WB����7�1ci��C}����G�rF0�;<�N?Xp�����}*��[�����l��O�ƶ�4p?45�?��ڒ��1��������*����؛�ۍs�"p�vb�R´'��V!�P�ӈ���K���Z�e�I�ƀ\�1d�J��,r�v\�Ys�f�l��Λ��T��'�Vioe��|t	#�h�}@%=��F���ɮ�=�n慚����^o�]��O��B�z�+ �\�\P�!�r�
�W]�
a{2m\��p>��V�����%F�W�0����z8O�����88��i��\`��\�Ǫ�A���I�w5���h5���v���d�>�XQ�pC��>��Ki���w�<��g��� �ʫj��O�6��۝)�xvN�R���3'_;�_.��?9��z��QC�m^���a��i��^���*�?S�
�pjT5�Js���{E��@�������fM�{K�|�ؖ�I�D�O����
&�Y$
����_r�<�SM���xy�SK�J����G��"�'g�^_#�U�*h#� ��ke�ǇQL��M���>����]��;f�^'YA�y	�c6����d�C&P��魔��ؚ�K�>#)A��|M�o8Y�jO���u�T����eZ�(����J9J�Ɠ�;:�f,C����.LU�Ek�����x�W����H������]��Դk�T衴��tp��5�ʓҴ�y�}�m�$��V�n,FJ��~VQY��'��`#�� �j�Sa`vt��{'�0����:>��+��UQ��RC�c���;2_Ŭ�P]����I�cAKD��K�7��+J,w��.�T9�h[1 w7��|8 e���=����P;�D��.r_?��0{,��^��k�o�t�3*��>�׬�ѩ(���\}�(��3!���^�s�j~�p(N̍�9H���;�>�� ��b�Ap[��!n�����wmt�_���y������Gn��3@���񥾝�����R0����u��P��W	H���?�/�O��W�xLe�;�30w\�A�?b�Ѷ<����R�����(E"�Mb�/���a��Y�$�G��u���g[�M�RL�3�^Δ?�I��!�{�/�Se����-r_E~ZDf��P��c�r�8NP�Nu��?HB�o�-�R�H�ul>lK5�%R��YKix�e�葒�#�踊��-�H�$!|�M_P!�W�G��V!���NF��w���36aI27�7Y7�x�3D�?��+\����nW=�+���q�������z��>U��=q��O"'���~9Ѷf{g�8S�`-�K��1/u\]��%����3w\�{�&;	Tb2ڐ*s�Y����'K���-uDV�x6r�A=�gP�c��r���	(�a���:,9�4̮<ܰr	��,�Q���$I+hq�Ǌ,6XR_e��B�6�+}�~�c��� B���܇'tq��]�8u����J�	u��'�2�}����źi� ��ɵ�~�2�WLFN��-	NMT�5#G�a{��,(�|O���U�{�I�b����uy91VT�=.*�$��oRspw��9��������k׃��:{�!]B��c_q��ro���M��	F{�#.�bs,��[���i4Fr�-H����ņ��|~V�aו�@m8#��/��q3����mf|O�jJ΅�W��3T�EKnW�Ш�js�9�W0Y��> �KCP4��]��/�NǶ�+A�:1�{�M�w������[L����0��sT�kJ�v&1o��[�n��*�]�����[��L5����@�����4e��wX`O�K+_9BI3��H6���8[�_1N3}G �a^��]<���r������QoL̰��Wm�Q���KI
�N]&�m�a�E�M�ۦ!y��2�r�@	,���JGGP���U�`�ͦ��ʤy���G ����<9����l�mH-M�]d�^��}N$p`r��%<>5L]~U3j?�5oC�"�'̟���{V�mC�}��7c��U�:�a��_퓪�ӳo�9����R`hH�*���s��k�א�,�Zu�~��:�va�.� �<�Nn8_�pg~���C���	�����/��9y��q���F�m��8wпi���b��-6
��wB|���@�$�S����t(�M1&M6�r����Q�Nn��`VT*u5X�ؑntO(��߼���l �|��)�� ��ѓ�z�AtI� #�X��=�S c���4e��R2m��ܷ}`z8�Ŋ�Y,c��~�Y�{�1%X�;���σ�N`�M-���gN��������Ń(�_D�-�SZ�@�M@�>k�Z{	n�ֺ� ����d��>9�{ˎ���_�<��y��������[\U<�nD�Vk_���KGe
Ц�1b|t�@9.#�]?����W)� 2.',.�+����ȵq�/�F�$xmkH
����`��"�� cF̲�",��L_w�
���L�k��U���=(�S�a��
?���� ��8��.Q��j�J���
�Iq�9%u��)�^���/�k���xn�u�H�<��w ��f��K�"-B�j1���]�'�4�9YQ�����~���)�00v�VJ���,��L<�[w��o�[n�i���.W�B�qC�^��ɯ�ΞY���t�E��˰�8?�/�?����r=Z�<��� *��'�~��3���,Pa^Ҍ�xЮ��1:����m���/��