��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����Q�&�$G��Fs���K�+������;V�P���l��X�g�rNR�;hVC��D}�LX���J�lq@Á]��d��择+I@��g�&�Nj�{q��"H_X�&Gbr��[��.$m� ������bO�J��jh�x�#GC��PN�����{"<�N3N�)�	˿�`>�q�&:Q �#�;��'b`_�{��W`�
jM��,�BD�@�pـl񦦵-Nz�c��.�W�G�I�p��*��_��
P���h��W���h���4a���gT������?�TB��\e�'��5b�D�?����@3�}P �H����Ŭ�#���V��U�J�&���)��j�-j*��t#Ȝ��G�՗���/��e�w�M>�� ǣ����QuОd�Z���C��|k�ů�$�|�͏)��ŌH�:�+.�O������wE8ɐ:N���\�bSI
s�C	e��T��`��#Qh�'��q�E<����w��������\�����;"�:}����������3&��2�64q;�z �h�!k���|/g��kʌH��GR�_���CU���8!g�;�t�����|E��'X�U�û�#��K�fOݖf�9���)��?k��<]�_��˧W��bGX��(��|<�D��m�]AO:�qZ��cИ�}�T3a��@6����1ۛEk&�*��cGerW8b���j�j̛3����\Ӥ	T4�2����|/�e��>Xg�B?�mi���"�s4��/1;Q�6m��˸�@"SR��A��Z�I�w�x:�u��\�s���<��l�mpϥ��	�<-��J
) ���զT��'���i��@{
)��'k�`���o��x\���V���̟�{ӕ�l���U{|���ʳ�Qt������Kx���SCUl�֚�V&�n�O����(1N���Z���p��qd�q��IW��	ߊ.e��`�N����C.�]TT��W|��`��i ��>��h/f������KCկ�~�>����� U�Dո�U��R�'�Y�&�N��y.Ĺ�*D��:����̄a�R�~�I�ΝP\����e��a��S��|L�=��B�#��%$ �u ��`�c��	%����&��{WI`x��G!�Z�k��@%+5��8P���[T��	͑�h�$"�\�1j������-�� ��V��������10B>�
!����n����ٙBB�N��"ۺQ%[C�l�SX�Mpi�l?�e��� �.�9�3�Fr5���=3��؞�i!30�޽��(���1�uƁA�pL��F��LNG�m?[=n��b�L6V�j�O�N�A弪� "�5Wg��m6
�?%���5}��7a4_�b���fx�%�8���M�y#� �C� �J�*f�b��56���r5z_�q\e�A󏕅S,%�Ƅ�F�_c���R��.L�5�~���9�=�4�r'3�럠D�)C�d�;In�K��'1
�h������ѧ��95e�y@��nPu�<�^%��%�|0��3�ә���4HD���	<�?�,����A�z� 35u=�lR��D^�D�|�F�\{�i LY��TEg�_�dk����z�ɜI���A�����V�\�V��C����ĥx<�9�q̗���H�l���I9a�w@U�R�
=���
��tz%�i�ژ.����~�0�IP�}-%�̪�^J�ѰZ��3@g~tp�%���2?�d�AmDY�22>ZHt�����XǍ���̳�gC��.�*F.1ƃ1�eu*M܊zO>/�J����P�X>����tᕅ��n*��˂���}Mt`8��x�+�f�ަ��01�Xh��Dw�Nۭ�i�����3�8�V��'���)S��U���Q|�,�����xf�$�m/nt]�Op��-:�X$K��Eć1�Y����ͭʖ����Inժ²tcw~:|n�T>�9Փ�Ə檩�}�Uv�ߑ���.�<H�i7$*:CZ=�?q�Y��8R����*���_�-%��O	�r�bV3��-oz�;+�JU�y����
ݴ��b{�,��΁^��I��M����6,��F����M�kuږZʆU]����EZ=6@hj��ǁN5=�iQf��̻�Fl�����<���5���E�c���+[�&sLh�T�S���pg$L2�{(��X�m�n:#�`�ld�����r�wVW+'rK {��nQ�}�i6����@��q�	H�
bލ�1�0d�
�e�6���Ħ�-T�˾vu�gA�uo�hDt5�J?%ۮa�Z�)�fj�|V�FW۹}�d����F�%��T���n�+S�􍸀���)�8�����'�����҇c#�պ���Ɣ���Q@�V��bő�?٨Jĵ������2�dD��Ѝ��Z}�=D����;�ص-M�[ht��6��=(��p��K���Ds�z/3P�2 L�7��]9ðSg��rv�w��k V�=��S~4$~5,H�J��i�P�I0�	D���6�	�%]��"@�h�N�B���X�8-P
:�J[�W_!�2/��İ������_dA����C�_9Ԙ9�S����e� �MB%��2-GEI�M��*eWV~�����b�9^
Q��x�y���P�)���5�j�(�5q:'�׈�ާ�D��&`Bn5R��Dym���&�
k�1�&������2 }�8���(��r�j�)V�.6o"ܾ]�b7��\B�}1."`D3��ה�ݪ |��Ab	�V�UC�?,+���BKڔ�G��*��7��p5:aK���i�|	!��	�a��H�l xKl�1���x(��ȯ��2ۗ3+�lh/N5���ꗹ���K̈�{v�4$�x��l��o \����|'����V~3�凔39#��%]�7���=�L)3���	���ܨ��	��qF���7X"���bK�eqq��BJ�f|��@d^:t��)�7��N���[n�x� �oR�20���k\�7��(ܑ�;�5/|>������]+��ѹ��s.�.�9���o�Yq�{�Rm��@�w�1����w{���qӰ*��1ddCE��{5�y�&h��g�9[���"����+� �Ə���������E9�mc�nqgp�=*�|�]�﹍�h����P�G�4KKjrg����'�2�N;���8{��a=������.�͠� �˸ihm@�B�Wq�6�6)�bA�Zګ���v k�Zѻ�����t3j4<��}����^= �S�1c?�!d�\j��S G��F�Z���Bip5�_E���ď���skH�*�%o'�����.?�;�7�ʙzy=��uߒ�������k�A�;ֻ�& '��	'��5�����L�OE�G��ҭ�	I&�&:��r��0T8��4���G���{)��T_
[7��*J�lSpR�44jM�^���M���]�������!of���ոF�;�f^t�����Cl���&�B��W#��AqC�d/^&�|�3�Q{�Bpu'�H
�~�^6���z�_w|�����A�
�A��� B@I(T^��FIm�����5��LT��q�n�y<���	g�30����;)xǔ�ǹ'j �+��x	Y�@I���m��i�@o�E�̉�8 ��99ζ�����(9��BG&���:f��@���s��/�}p�Ċ��!/�n4�Z�I�R/2�ԉ\rQ?���#��ȡ��X(k;�S�R��	u]��b�e�vLjfA���CK�j�+���]Eͧ��� �*|�G�0�@VD%>ׂ�/�K�^R���c���I�`k�����g�Cd��B���=W�;)�J}s��μm42�%&V�D���UQ�a�7U]����Ѧ4͌��R�]k\��Pk�1(yT+3{o	[:��x�`�xh F�<���lL�����!^� )+�7F�-Ӊ݆ٹ��Q	l	yx.@X���k��U������W����/?����Ug�BC���Ųɢ��^ќ�����~��-�w|�T UP[.URtv�p�ĥ�7p�4��'Sx�!z��h�n˚�z����i?�&��h�(��q�:�(_f���;W�sU8<���
��N���T���毘1��+�f;D��~���>�qˢ�Vj�K��R�����0���������k����RX�+����4��#�nO�q%�=��	-���*c�ƅ�ȮH��ڃZh�O�	��� ��L˰�6|d�P�aE�E��"8�P���֋p�-�Tϛ�#̄��->��<�ih-��)�m�;ff�ͤ����);�$����i��@,;i4���+��o�E��ݡCE��L��}��PU������=� m���q�5�h5]��5V&O�MBN��+�� b�+�gjI���	����0�q����S����>��}J����۹�U������e�2��n����:}e~W��1�"���4|�Z5N�:Ɗ	�l;���M8��M��obA3b�U��|@|�*{�W�Gcx�G�Q�Fy���u�([�F�g1�3s���ϋ�/'��y�4ұ�}��D���<�ab���-��$$l�q�e6��$�p�����(�/��l+4/Ej0ʷ�hЂ�D� ĉ2oζ�?~����2��!�u�Y<AL��b*�}�	:W4G��ʝ�?���	�0���F�^d��tꙖ@���'�5�hn��'����wMns#� �8i:@�@��A7�e�E=�/�,��a�>����JT��ݯB"r��F|�_+R���.y��'�v����B���X���C�] �\ݵ�@Qm&0���H�d`OR��Q����s��et�������N_|�Ӽ |�2�s��x��b`/E��ܮfꓚi��������RWZ�m�;;=��qT�Fi�'�b�>U�f&�e-�kK�"�W7~!V*��?t�r���Q�Ϧ{;�j�z�i�x��d�&��~𨋙��Z$ǫ�K�́��{�i�~����_lP�8����|�DvIA��m^��W�n�g�[��6�7��GS@Vg������ޕ�%J"B5N�]�^�o��=a�1Ӥ� Yb�k;,6�U1�h*��� &I�� _�j�^؁S���Պքw	���\�����
�ȏ���S}%ǛoX�@�Z����=�Ncџ:}s2^��Ob�8M�M�NU\Y^KY�3����W����6�g�S���_�s�)�V��EOS�����Y�$D�&����]y��$�U#����3v�M�)���(��e+a�-w��2RVO�����k�R<�HR��5U���|?��Ğ8�gi�l���ЊR�L�~tiU�Kg�%p!�=n�h:B���@�Ά[�|��u��<��P��W�l��I⿈��}p�݃�/��g�
8ӸQ!K�1d�R������Ⱦ��
�;"�h�VZZ�8~Ĵg��1�xWB���l9�S�[$�а�Y_�w�(S���,��r��~�x�V�L�� ����W�F�?��y���GX��߿4��
��O�������u�OZ�pBa{�/Q=6>���}!�W�,����o\V�� C��hL�����n�LrP���}��5�����z���?��7�q�)�G͚ݮm��'��N���D���>O.L�?�!y78^J�nFl�XE�Zb�y:N�xM=~�ʧ���t�K~[Q�yf\z Q��~v��tb|d�[&\��2�
�wl���IT]� �,�5�M����]�b��^���y�{�#ӻV�x���O�����BiX����F�վ=3�c���( U������L��n&�Mj>J��(��^Ӎ$J�-^�ك�ݚ��`��D�D�/��7�,���}1��Ў"�1ӥ�C!!j*��-�� ���ϐ�������NDc�'0�R���$��8��?1�&�����F6�A��6�w���Ӛ���m;k6���*�%F(H�������s���H�K���w�tg���o�F>Ţa:�Pf���Rw>}8��k0���B���cb��U�INm�\*�s��=��2q�Q���̗�/8)�`H?m�a䙰�Lvr�aLE+����L$E|-���m�˩�D���ν���h�N��;2u'{1��1İ�RG�s�=g�m�"�����c��qk$I3+pRz	=W�䵊:��fuT����J��K�kOruU�ö@�+rC�8��?$	i����AA&`��P�k���R�O%ע�u9gDҺ�K�ƛִ�wQ�y�C���=t�]��@\�(_�JR�o��� +�X�<�N_]�]4�.�e ��g��,X{����~�Z��8��ɸ��)$�)�G��u��Y��c��N�0 �,L�nB�_h�z�z�߳��9?���jR�' #����k*Hv=K�j-��M4#1+[yRĥi�j�1��4D+"���FmGS��!$������l�m:w��\��Tr(S��'%����q�Я7t+v?��W�UR�ءE.0��y)98 o���͗��9:-��ѐ޻IXSR�N~��a��<��:-V��~�+*b�ˤF��QK��.�~ӊ�n�ce��l����_�ʈbQ%�PQ�EV�9�Y�(�o�@v3D�3�����EG���!oF|�Ӥ[���d��a/�nNU��,����Z��W���"�����SPr��sQ�����S����gxH6q�Y��TR����;a� ��9�z�{�/�3����>�,_��<�����b�\4Ӛ8$mP�b�+$��[pI1i��?���JΩ������%:X	�ݚ)�.ь��;3�T���_ʾ@YO�BЩ��l�8)�hƒ��@������T1�z����oG�``
#��y�$�Yֿ�R�y�������ʨ6K�bT���E��T�^u*'��co���%wS�A����[��������l�i.�H�v,���{��Ǐ� Ys��.#��ڄ�L�Y˧�n������&���8Eʩ���>�w�9�r�t쵀-��KK�������x�������;ϼ�8���[������A�[Ӫ�d���t3�1-Ȯ�:��];g��H>f��q����0�hUF�E�%�JO6콬�a�~U��_3�.m
@�r@�����nV���񽇬�2<�%�Ť��I���L1W����̅�Bl�v$��l\�O�
�&�n=�d�:G�T�9>�r��u��Yf^��ݵ@�D�(�B?�'���:�l�It�L��S�������7�N,�ťߡ��~`�4�Q� ���ڤs.�����C+%q�D�0���m<_��Jtw�	9�L#�,s �K��	�]&�=8�vFDaq=d��(e!��ݙ��T��4{�Vb�k�]��kt��lA�	��M���	9�b�W��7	7Z��m)�@8���:�#PƳ�}V����S���TQ�����������)��q[1�6r���j�>�ݛ����AΜe�R͙*��&�3�_S��O�'6$�1e�a{�.P�|������fba}�,y�	������r^&��uOR��5"�O���<z��Ro��"�2v���b'?]��\�!�(��,����/��Z3A�z~[�J[ձ�f9Af����=x���A��1�z[Kv����H�O� ��"��/l���d����@nk�k6A;W%�ۑ_�6�QQ�{��d��V[�m����\Q���2�+}�~�#G�#���Bk��I>��F�6�s�"�ZK#5���kx��-�{�?�0�
WvX��X;h�G�	 �����3�;�
�?���V��*N�x��Q�(P��!�l��Hf[ ���PԆ�W��p���h�+�LaRxT���h2dB>�p��I)<��0+%=H�5���R��CI:h0���+�^3�Ļ9�\�̫�v�u]k4:f֖�s����o�X�L��x%�Y6�;� ʲ�p�L�6�zm��;7���ڰ���yd3�����o�_�'s��y91�P,^U�z��8@�E[��Nu;�F�%�c
�ގ()2��ds�0�+��A�@=�.T��qm��7ei��n>w�4~Q�>N���tfx��E���m�	�_��g��>O�Ǿ�|��/qm��HBP�]J�7*�`�`��*\��TNe���`#n~2�k��x�(�@�s$jT�q[.�P7��Q�{�kU% x�
0�Dp��0\�Qm9�[�>|�"����}!fo�#9�g\�>�K�'�Vo;�{��+�xׅ�ږ#Xᇤ���s��
��������E�ϑK����p���+Ԛ�$)��5,5�Y&!�#0�*|��EI�'f-�D#}ƿ���xj��FI.גw�P?�l�l�ê���\P�7a<h(���]3�\����>�h 8|�$�V+<�����M����+O9xɫ��/ &&�غ�g�4n=�V�&��z8 �o�P��ت�s�nD9�B�s�ޖ�S��L�8sֆ��a�u8'�]�y\^D�pxy�Zp�:p�zг��w���~Rp+rn��6W��B�H�Yӭ�4CL��KM�4�v�s��5~k\�}�&�6�0>���G����������;��,["�Mȳk�*�f�ǻ�����Pܽ���EK�u� /P��ɹ��V��쯐�_�mj��c`����*�=+�w��� �Nh"s�?K'�W�m{c����=�P���Ss���&�Q�h�
��w#>��AOrƭd|������������܏�mp=:d����C��H+����"�8d�pèd+va@;g|,m�Z38����`	��ʽ�DUNMX@�n��+0@�M|��tő�f���?�]�.�ă�@(o0�� ��^������%�����G��s�yn<�&��ﭚ	ڊƏ�N�r��_x������D7l�,3@wb�X�,�D޵W��t�Q���֞=s�����-�2w�?�'��y-N�%�A~�&���=��fbO�^Hň��W+�Z�;�6t�P���A�z�C�j;���"�R��_I6?ZW)����w䐧55B˯�i�2i�=��T��D�U��%I[H���?e�q�c_th���H����|:��&$Ҝ��o�l:��d(1Yp��"�Vg/�&�#����/�u2���-��t��Gw��n�@D+B�m�����??��G]��/��fJ&0���=��p�=�S1��80�+J�;D�$�nL�����͏F�q�R�l����w���t�/�P3�\%|G"����w�����f���k�}\<�i��hfr��jC��%O)p���� �y�z:���85�8�� �h��R���}��+?mi�b�"} K�y�8��;gu��lv��,�M<2�>9&� �e���Y�і������]�;黎��_�7h�]w��ix��xWnt�A3h�,��r�#��ۨ�� ����puճ�r��ˀ?������=��/�0���.��iSѯ��A�gF�Siܶ�)��r_�۝i|��ߑ+����8�k��;�&�IO�װ�Z�N�&�gǡ��ct�T�$��sv@W8��k2��A�-����~�	�X;�p@g$Qs�R�`�RYm��\	����0ҧ��p��I���+��8PT�TF0�`-�2�2:�jx��5���f΀���i�l�\.w�����������Om�������<�iJ�R|��.z�rvZ��;�9+��榱UE�/X���1�H����fՐ���79Z5Q�|��ٙ���>�@��6�������YrĎ����:!�s��D��_-��`��ѷ��ܽ;/E$>Z�%�D��Z
�ɥR��Z�ԉ<L�e�w+��`�f�j'C��\��!�S�Wx��_�'j�׶�������<W�ЈvGZ�A��'ƵpSE�	�h�ܲ*z�� i��l��[ݭEXdm3*XyϚ��v1��5()2l:֩���{�h�w��*�����?���nc�j�T~ �g�sxx����n��}��L2j�z��^�a��/Ǉ��_�������B?2F��nM��w4f<��m����e
l���H�>�-?�l?�T܄��+^6� ��Nn���tƩ�K��뗶:�����;�ī_�;�(p�͗�F���o���}F�>zZY��'�yQ��P��5W�����C{�3��DIM2?��V�p�#��4�˗9��7�����-�y���e
�Y;��l�,��w�>�P� D`\
������x�Q��O~�z,�n!�D���#���"�r^X�1���:���{��1�+ ��w�:�eO`��K��if��B���u�TU�s��� �C�?�M��f��F�?�-�L<⯻�zsi,��W�%cć�r����$v����Pǖ��2�샹 ��T�����J�U��+UM6"$�ϲ	N�!���G�o����>��i�'��npMڙ(�q�ғd��ܥd����A`2W|F�!���}��%�|��փ�,�2YJ���@��>]QE����a��]T{��'�֐oʪx�o�мJFB���Y; A�%���؄.C��j�u�FX�t!>��t���k������Ǥٺ�)\��1���O�Pv �/���5�ו�������z鳾=�@��wi�|�΃�L��@~�Y�8Q<P���3j\�d��*>&w����V��m���vy݃��>��l�Ӈ"�TwN�W8�*/k�]J���Y��!���5M^��N�=���t���G'��(zd>�	B�0\����'��N���r�)���������=�׃[��v�]t*��=�M���JrMߣ}��9��	Kj͕>;U\��Ȫ�[�9����V#f_�;�]��~����y��m�je��6X�0SH0�ۈ#XM��W��>�?y�8s^�ۅ��z��ğ���+�T�m��b~�q橡��t�Wr�%�0���O��r�uI�!�HF�,��>�\u�����>���9D�Y&�h9u���J������q�N��ywwp>�t1:I5�nO�@⾶J#"f��0RtN0eg� ���"�5CgjEQ�:�J��Q��Z�Wds�JfPz���1��s`�6Խ������+M��y�ɽ1�a~~p�a�վ�,^���0M����h
f�@Ղ��K6�ܺ6o�q��g���rL1bZ�|�LF:�QE�?Q8��6_�s�iC&~l�v-U߽��W�5ZH,���Y��y3�>��C�]�S-�K8l5����ŇOී���\L�`LD��j��q$��d野}�����D�x܌�����&�?�,V/��y_w��6��-�����b�x&�lja%��}�� �����V*�+"[1fb��G��^H-+�n������0o��Xf�(U5f�1���~�\�`��
I�r@��u+�k�=cs�k�R�4��z�d%%��^GÝ����C�o�Z�oh@t �Z�*�
���.��ņS�3�(K)[�&s֑3ݝg������F��S�6�P�'���G"-
N���7�����\����P�4,ވn�ߔaQ���F�@����0]�S��2�╾MI�#K�B�e�$����:ͤ�J,w���D�NT�r~��]r S`�����os.�\O�� 7+VW��0�ؑ�ʭ�@�~��ވ��z}0�x��l��1�
=xtAR�7g,��H;��=&��I�;��P��q��`O"	.Q8�Lh�Q@��
�����q��6h�OX6l'{��G��:1�E��5D?t��)t����[����XX�s8�����*�t����#M̨n��s8V��"9oXh���@\?���z�p~~���l}@���i�F-��}�o�@�h���o�B6Bp��ذ�t�KJq��Q�t�K�\�ۓ7�Y���`RI]���0�|m�ص0��'V��ׇ��e��a�+��(^u�q�Yk�����Ŝ'����SX�݇��ez����[�(9ǔG*�Tw�)U�tgZ�M��[M{nyt1��eܔ���\�@ˊ��'�`��4�>�A�/h�,�5��n5�M~�V��Ǽ:g֪ݍ��%�n)��������r���1Y�,z�kSͣ.���-�<q<,���.q����j7_u��j�C)Ԏ%�[x�u	
)�>55K)��\4b(��������3؀5(5L����K;�ҔL�>�c�!Җ�[�w P�|����rѹ�c~o��@���zjb��ϞL�����`�JyܠMM�͢�-P05�4"6aDS%e�>��L�̼�d��3��p(�_ǃ�*C!��C�6��q܆s�*���)뭈����	���s��S���1Y+�N�S��}�T���`$���F���T����g�Wy�2�|�'����(� ��[ �M,����d��EOk�����0p_A�Kky��M��@��'Wk#XRR���h����x"y�=pӞDT	�@P"9qi�?���@qf�d�o�V�$e�c}�(��Y�pg��S�y��~,l�.�*x�1��T�$A@YЫ%����`D.���s��\i*`�[��c�ΨAi��� '.�7�Hb�c���V��k0�{���[ ��+�������}`T#&W|�B1�jW�/!5��-V%�	'��F����
��Zl�ؕ"X���/���Uh*�J0�6��N� �4z���W�q]	�Ζ*�y�_�2F��K�Cі�1Z��,ϔ�N��u1�y�>��E��A��	ZhD<�ɷE�ʙe�G��+cL����<���?�
���}v�-D�a|���xLC�C�7��ݔ�������V]�������.b>xЂ�l�ݔ6D&����H������C)ؗj��
6��t+m-���wxyy��*�{�t��)H��b
��LnJ4���d� �8K�wL�]�����H��X1P T�t�4Q袰AZ&v��Hn)��P��k�C�~'<�9:�t���C��0��	R�H�!��J5sս���2H؆��]�_���(�f��ZYiW� ���@�ʌ���t���TU�i���Uߠqk�;pub<��U��	�-�s��/+a���.0�=��A���o-lm3�)4�o��U[��ߠ�1V�	!E�yu�����ȵ��+�k��dK<I�_��������U������� ���N�S���w��/���z!\��Q��Ԫ�1�*�1Š.���_{*��q6q��_]�2����Xm��oEY�?:H�z�4����eP�-Z$��94q>_�+�I
��)���P>Ho��C� oO$���2Ke��.G����M-Z1��2�p�a�1�v�`ݻ�I���צ�A��e�.�V�Z��r@8�'@,;jg���^�����A(_�.�{Y�5�-\w���H`�)�:�hD�]����.�D�w �?�L����v�\,`���km���H�jL��YWB�7lU��,a)0v��7^.ƽJ�|����4���NY�a��,[��Ww�U��m�(R뚳��c�nm�љ�����O= �@�e�7X��Swy����O:\�����/�H�dmp\a�7��J���B+gZ�|ҿ��omVo"�2K��O�%^$��ٗ��������<�Vp*��y�������yO���zp,J��
im�T���.S�l�Nr��[=zI�~6S%7�jaZ��|ӎ���N��+�.?��h�~%�g�75�*9��:�ں��5��Tu)R�[�!A>q��ꀗ:ͽz�-q�ʯ�yt������*ȇ^f�\�8O����Yh*�����
+�\�w��;��5�D订���ȃe�.�j�]�c��cQf�M�P��e��3�{�>Ԕ�q�vB��V�'��y�	)����� k��Fdr��D-�j&#(��~�Vi�tB��i-sn���[�*4P��5hFYz߼7�-c�؆c|	�l]�g7��UK�U�f�>�n=�vb���n��u:�_=w̖}�z~G���tx�m�V{�ָ'7G���E��Ȭ7���|��?.�v_��t�Rc�43���>�'U��&d���RnW_���ړq���J���R��j+�!���T!K���5Ŀ`=�AHG�] �z���_�!��<[�I� �n+G��m��U? �IU�ͱ��s����J8�#�x�)Em����˨Gppy7��fO�߀j��xr�m';H�5�p�\�19�{�%
R_�1(f	�á�7u���t�}e���R}��i=�
�C���(f��N�u��Y�Y9��b�c ��ĢZ2��/�HU�B�aq�e�I�F�\<W=�h-I�m���!�8m�æ܍x�Cܲ�(H_�X6V�Զ�����d]g�xx�ԼH)�~ᛤ@cA�?@3 ^ �$K��iK��x��U
���Wֱ.V�'�Wܱ\���<zG֎/�%�!�{�y� ��a�~:fS���ئ*��x���# ���!�$Q�
�����In���D͏�JC��^b"&�'Z+!�
�<Vl7Z�_O�!S��lU��K�Deߣ]�����hn�,oG�bxkʄ"�K�����1�iD$UP�
~j)�%o����EC�]�ZQ썔�aQ�����x&��Zd&O�|`����k@̑9EC�s�ֵd:���5��%�;�=c�5N5��Q�#V�Ɏ��J=��G��;r��dDw���������
�fV$�-�j=�o8�D���*���U��7��=��m�]^v�z(v򈱲����ە��P��`*d� -���M��4��xIh=�ߚ̶E��B���A ���f�١;׏Lo�-/OR�\��_&��t����l>�e}�F%N���Gh���K%*�PU���[���nqqob��ݏ%��G�8ڃ+{+r�����r��,)�������K-qF��&�̐rr�7K
�� �h�%D�b2������Z���_�$&�T�<����y��#p�I�,�F�3���1���1U߅Hh=� ֔�*vJ��>o��;����`D0N%���]�Z$�����M�J��K��v!��C��l͇����z������x�f��O}��/�X�Mp��i�Jh�3�w�ۙ��W�7ti��m�3�/_֙G�R�T���	8:�^��!e�J�����a?��.���/�B2�g�ʾ��V��>���?�/���sm*0/㗳1;������T6��1$S�3h�O���E���;	!�.���h��Y+��?�%L8�HR�!*@f/�4�#x
_3
r������p����mI���୔�/�|k�+-�����S-X�*�m�Ie���gzY䱋=W��8��7����*^:^�90��Օ\�9�&�^���U@F���5,����|<�����hZ���Z� Hm瘄/�,uS����-S�g���)��+isc�3i��+2����'���׵Sv�X*Ǔ�`�NIa�����ߕƁ��wk����u�v�@� ��X
�y�Au:_U3���^dAnuFJ��#;��E�ל u��'&|���gة|�N
���4�b���BL~���m��*'�$1D��j~[e����
��']�i6�0�&��L_ڦܳuu+�T��kȒ=�a�tK��{���(a5�ưT��T\��W�����Ϯ�u��	��Qf���M<L�P�o�� ����v���A�[����!�;	�MR㪿E��|%���K�9t'g.�^_S��~R�
�hH�
�`�u5x,d�l�x��x%�����ɇ�	�ϲ�S��>�F[��z�벿��y�\�C,i��ĸgK�s�xR�II��}��`��MF��eI�+u+m���`�F�;���hō_�K4o{�nH�A%kN�ƫ��؎
mN���	�6t[�	���<q����[щ�>�hW�%�,�Ά~Ls����}����K�����di��I`�|��UP�f��2^h����Vu �I�V:9��/0�H����m�s��t�a�|��-t��{K�ݦ�����{���m��.��ݣ���;ʀ���t�Z��~�p���`����$'��5���#*Yׄ��G�Ŝ��H����=y�M�$&�C�	��꾫x�	l�0�r�$S��@F.��2�>���� c��a
5�(�y��f�LY�%#Ǘ8��@y;��<=|��V���Bv�M!J�������1��ÆOe��r�̟�#qƸ6�p|�$;����OK ���lK�p�b;;��5�E��H�����D�w�#f��l��u�q�/*���m�l���]�����G(r"�2,ص���Ԁm�HR�C��4b&F��눒5�*+GV��?���SƇ��CN�v
���:p���`=?��y��mq��J��k�@�wؐR�"�{�݂��ET�ؗRP�Q6}�l*�ƒ�U�&z�D��=��U������޺������g�w�l�)^���ŉ1�.��*4Lô߾�uӞ�.,!�Ӳ4Z46�Bv��1&*�3.���+h�4c�Mlg�O���u ��d��¶{��O���Q<Q� 02����1Y���3�?"̘��&o�Q=RLv��$^~m�/�F�D���D����(���R�ӡ�G8�f���s�SQڲJ�!�x��D;�1�:�ӭ��k�e"KC��_T�����y4��DOvv
�;���_Ե��Y=�A��%m�+8Yt����qKt��d������5�͢+��8D��6����&?��?BZ��50����1�؄?�J�\rh��Z'oV1���Io�K,O�n�P�P�@�� F��X/1�*]�bUv.��1���Y�77�W��)�G���3%c8`�Gpc,�H� Q@s&�[n���֮��k���R18Z�w����g�rIT�[����^��ء~I�m�ծ� 5@hMN v{8 BiecX�߉���ey��ܭ$�WzȐͯ�����%�D��u
6,�z�1I�7�:\H�2�]fd|�6�ރQ?�uٟ��DH��ה�՛��Y��k���:��`r໗�J�&I��GA,Ln����@�E��:
�C�&{a�����Oɛ~��h/M���4��D���d��a9�t�Z�Q�y�:秲��K-�i��cc���?*P?���6�%(������{lsvNW�����~�/�Q*R�	JɈ�O)Xi�Ð�uX���E.�<�.L�_y�˳��F���4X�9�ct��̩�:XZ�L����(V�.����0� �s ���*������vC��n$�ja&��;���7��v���ݛ+���'�
�}]������r��\X�P"�����,<r`��c���i�#=��l��Aw^�+&��
Ю� ȶ�H%��_�ݑ1y������\]$D��У���]�E�S^Yi�(�g�mG�=\�˳��Z���.-p��bd�`����t3~pX����2���k�UM����5���=�Y,u�λjhЌ�@_V[�|�����Z�nt��b�@W#�"�T^Abz̢��
�]��eF'G@�{.��{�3��պ1v;m*6(D��5�E�x���3>G�� ͏���biy
Q�i��!(�Uk�"�*m��04�$G���F�k��5w�l<�M,4��sAz�	Q����|/��\ۊ��Q���䤱P)P:�`��0FWN8x c�&��j��6Z�)��L�솀σ�}���t+��h��b#jV,2�D��Sl��g���Iʓ0���!_����I䮧�)Xͨ%y��$&�H�K���/(q����3�|o��p:��T�]�� g2=�RR�չ���c��%2�go����T~$TW��(��S����YX_��!Y�V��L�����{0]��O�k�2U����ڍ�`�s�++�BDf �-��
���`YD��BQ����yl˵ܟ����oT<�u߷,��8����|Ņ�^��tpI�����1O��[��z�����	���s,Y�
־|�Pr� �gcL�s�\q��G�x��I�,g)�<��>��>����U��y��!�"Ix5Yhv۲u��]p	\�Hw{�Ν�q�Ne:I�H)K����,P�)z�CsQl�so��%T�=�\���e�LC�ӝ���<c����ŕ�R,��@Kb�E��aג8��>�6�)H��i���+�p�������D��K_���,�ۇ-)���'u��c@в�����[�w�'��J~�_�p;���ϦW|����sPQ�@��3�O�\�-�^�QMvy���yi=��xHp�3���6Y`��4�n�+,�8zu��$ �f�7�g�(h���v��D1�~���߉.2e�%P{��W�1 D��|G4��h��:S�^�i�8l�^�+ZpKU�G�z�X01621U�/�쌙�������>��̫a
�ц%.���C5���B�2(�lR���Ҽ}i�k� ��n�bN��*j���0�Ҋx;�lF���JWi
oYz���0�`
�I9]�O�m/�[�}�7�"c��I����jo�����vg-�5v[VS߿�*�g�K���w�=��4���M�3o�^i^���.��8��n�ř��0��O(2�3�,����"О���|\m-S�?���3V?�}���y~e֔pm2��3`�U�Kh�i�*�fE~Q<;�I��z�ё4|^;qv�+4X�*n�ʻ3&h��wSX>�`�ц�� � KIP�@�.R#,�L�X8��e���[���(@3� od$ެP��(��Ib�i@l0ܵ{��T,{�ž՛F�aD]���Z�f�USq����^����c3T���e �$�2L��='�D��f�$�`"�Y��Z�dQ:����!߿|�F���Ĉx$����V#�T�x��pGjdY��Ļ�X{�(P�F(�lP���o�з�g��g�'2l�T�ahn�^�>;�+��L�
	�F΅z�rZ���U�`1D��hH�����[.��ЭO�f��8%U?�H���ǐ���ο���^�����w"�T���g�[H�ޔ��ӯ��~~�%�r5��:/ڥ�Q+��U='�|�	��`ֺ����߼���i��Ԧ�Wdl��u���<�GT�/Ҫ��#uŰj�L�K�ՑE�<�ѿy����ߏ� y�����_S?Q��!�-����N������q7��u�S�N,o�iQZH�+�/��8��'����䐾L��0x!�C��?u���m�9j/��i�������?�J*wW�A��T��e��͚�����8�<�����y_F��	?��E�5� bX�����R��$qj~���;˙���5E�U��\�їGO��D��M65�Uui}M�4Y�L1���yT�ZB{1♯��ԞI��7PC��]�ʹN���7�����	d�L�ԃ,`���k�ӗ�؟ 6Q�GHR��sO0��8l���f�����r^�@x�r���"j
�A�1�Yn(��5���*�G�$O�h����g�E�Q5�L��h��J���@R?s����í�5��ԝf�Y�G�M��h8�=uj�0X�|wJA�" ⺧Ä�� .��n=�ϑ�B��c�{�մ�0:Lѡ�{H�	m��XB���Z���p������{4�Fɋ���((�QrU�1�y�+[%��&��e�ؓ��k��T#0t�$J$�.<C'ז}h�)�AtZ��8��~_���Q%���k���(Y�FZ�B� ���З;v�K���(���l��:���E��Bۚ^! ��\�a�J/�Iͬ\��1l���]ց`[!��Q¦�4b~��/��N�)����cD/=m;�Ɏ�^�sσ��]_��r6�vT�N��^����ßp)�)��c�z��m0��<� ZfI~0jF�$�VV�.$5�M��4z���J�<빻"��������8�6��Y>]��]@�zѯ0`'P��|�CK�������|��LM�U?�̺v��H�A3/҄KO�Cꏞ�(�\��i�x����^2p�W�Y��d��2侜�(�¥�L�]�f��0�2�,��Zl��Bt��\dv8n%Z����BO���������p��V�%P�l.�l�$�<�}oc�!��K��6t�tH��;v�q~&Q%�{�}�{��|�ܘg5b���4��,
��nX�]���t_���I?V@����VmR�l�k<B�;:BC�!��{cG�)_�/��7��d�%G�щw�@)jH�������<ɹd�����?P��|�nˀ����k_�j䕕�dH�	gH���씈�7��40q���R�1�_c8�Ӟ�����[�{��U����K�ؒ��i��kB�8��S悈ߚ�i����*
I�x����xI��X��2P���i�46�l���E���p����k�6��)��������t�86q/+��`>;���:�t
=��j��Kt��m���@�lB��tʫ5�xM@�Ս����Jȯ�]t�sqv�r&�ʡ�U?vM�F��J����C0�ٜ�t�D��E�cG*����x��?�[B������a2���߷�o�! �²<�fFb�՘Gڇ�k/U�c�b�A �;��-�O�zhS�^-4aI��|K�pTI�'c.\���T�y��h���[b��=jÿ�pL�7�Ю�dph$,�x��mPb|��$�_�9��e�������� ݬ%b�+$Xz{
7��"�0�X�+ln��5��_��f2(��t�a;�5��~��e
�"A����X�r�4�h"}�	���n�[!d'�c#�����(�r�
n����pF�|i������X�ך��m,��ޛң���ۂ��0�Q��N�	� g����]?럼
0�Å@j�Cdæ�?r�5A����#���,��Ijæu��`�WlƉ��e�~MCO]��e�2�6P�t�@⤵:��Q��C�5���-Fu��¿�����q�QI��S����Qq&������s�Lr� J�2�y斡����H�h���Py.�m�|��c�p�o��=�"*B�ȶ�_)JZV+�؏!���T0+��� `� �1B��R��j1N�O:�pO�]�(�ryTţ�js���$��r�y5%UUIۼF�K
+��E^\�D�C+k7{�z��Z�+Z$���Ħ]c����[�#�B��g<���I�{�2[(�C��[DƆǒ��}�r�����o��Jt�oՆ%��;��,=�il��xKL��f�k]�� ipe��{�\Ψ�}�rs/wms�
i,���
	{��{�"f��cilh2E-B��#�'s91O�]&J��g�l>G/����,�N�������8�k�R�zطtF��R�c������Ȼ����b�E��ѻ��#����۞��,}J���4^�u�9�S�0#組=�Y����s]ԝ/
�7D������Q���i��g�bԢ�����X�3Ԡ�����M
>���l�\��P[[�&B<bi��Z������8=���=�Z)yѤgߥI����e��� �u���k����fz3�fZ��b�����O��+S������������f�*�w}�2v7��y�a1[���8�I@+�mf7�h�!��֠#IFQ��B��g$�pJ[�u���p_L{�&(g:�9�Q�M�� $ ��Bt�~^�},�����u~زN�<��F>0z���n���da*�r����/���؎�p���Q^��dg�g��}��
����V� u�0Þ�y�"ȹ� ��IIj}u���=�o��U\�-�Fa~A����ϵ�n��u��66e�J;�qf)��g��r�2��&�
���n/�(�;�����X���XWټ�x��
���[�J
��C�	��7����5�O:維s8����pϴ��T����p
��|픠��p�`�¾��Ґ��T��]#�w��,�vE"�������6��6�la��f�JCc�+,���Ø�C!�,�nGx�����ݵw ��1�C9/����st�{�L�/I�9U@���&�6\�)!����V%T�%N���5,"��uٓ��˅�o�Y�������D�T�5��� ���5�� /;�&b(_V��u+��nƅnڟ���-��R����G-�N��G�,�L�P�(ց�~�K�t�_WV��Y؎����2��ΣjN��V:��؏]�<�y����B֍FVr����z=��t���*�Lض�*_��3�d)к��7+�:|mb܆KK$����FW�x��T��|���1#��3��A�����d�S�cE�w�sLO(!�$�/x͍*���[��UBZ���
U�#^�e��iSRg��'u�P�x�;m�I{�؊cA�K��Xa]��#	�It���?o�Z�!��+1�'�0���Hr�[R��##6�&�XBK�\$�>wȄ�~UO��=�Jl�z
O �ӓ���3�Wژ�����Y�i(�.�D,s���?%���3]D�p�Y��Y��'��}� #C�F���TL�<��N�	�����Ēl�'Q��2�b:��R�DV;0n���9l�((�z����@֎q��f�G�ϻ��2�����P@�;�C����o�O����>~��m���.��ߵUW Q�~b/(+�]qZ�+ғ���GP&)W��a�����&�ʚS�'��¤'��3�?pX��mZdr8���+���JT����y�a���*��M�Կ�R���ݒ]e��I�/j�B�̓��[�H~٨
�ӛ�+;"{��8�{ ��؍,�����P�0�o]_�
�H�<���s�jE��y�:ma;b�����J<H��6"kj��!�.��S�3�ι�,̋Bc�P�����%�?A�dy�E�t�KLa4�hi�0b?���)�G��S	\�d�p)?�l���?{�b{�c���Ȩz�[{w��
?�A�X���|@w��Y�����j�릃����܄��%�8~_NMKeJ���ʳ&B������3����(��B�)7��t�l�K���z���a*G�#��󦕗!���ק���]I������D1����a����&�����Ӹ�(�3
���URe'�nO�d�{�8T(>GHWz��+H�:n�%X����\҇Q�I)troK�h�`�I��I�x�zP#�`��;�&�-������"(v�)���'��H;��;,Sz���W�����xx�}5��+�X���~�F�O�O2%����M��/�_4a��6�� �"��9`����
�I�*�ݶ�l~9�L��H�a�f&����S-�sjuf�%����w9�)ݑ�"�����/�|�>Z�H���9��r�b��'X>��_�6B�`��Z���,����(c�.�)Q��,S)�N�*.D�-��Pd��v�i!��;����Z����<뇏���D�����8{� �*L�J�N������ԙ���Χ�8P��i������Fea"��Ft$r�P���%�9��|-��b�R.!�ʹ��6��K6���|a��I��_���X��rm�iy��Kt�CŸ�0�z`'��<㲵m&Д_�i8�y+1v��M��m�z)�������V�1����:/�@a�)��ŊKV��� �J��ٓm��w���m��bo�>) �r6�=�<�*Z�ޚ%��oX�~����f�����YyG�"9���H�&��"���y+r8φr'�RϹ9�� ժ!�)�\C�8V���SH��S�*ZјKU�-Ʀ	������{Ks=��x�0�n��M�F�������h���qo-�w7�������-����-�b�\�<��ڢ(�cGo��yz2C�ۇ���E6C�}y��Cց��&��m��A��F,gMU!͊���@�ܐ7�嵵K֔N��,�M�VM?�k����`�J��'"����13�Nb�kv���U&ʀ^&|��;\�ױR�>�2?g�9D��58D2�Fw��$,1:���3�m�MI��a��v��ئi&>^1n�"{c����Y0�0���-�%>ѝ��~���p���Y|�u-W�KO �h!/g���h
\7*|WF�/�\����t.��������{����}����{�p�����`Y��-�5/�-�7� ���Uw����_�����X2?Ѳ�ZH3K܇�t�,�=�U֔�F�ڀ�b�����uM���_r0�EF���ԣ3�͘��ē*��!��)x�	������,�eq�[��C�ƠF}2��[�(JRn�����i8;�ׂK�sWj{��n�˙��>3�JH�������Q-��r����F�g��7�����<˸����Qr��n����|gh�\V=�y߫>Q�)�1P<D���yj�V���B������ۙ��3P�R�;3�+@\�U�8���l�
�@�*.�1�Rq�7�pO?��-l'�>��9�zI�3 ����Vh9�� � ��V[":a���}�Z�E��!�	 n�����9U����y�fV�d�����{2%~��|?~�T��g�������d4����hĮCM�Y�A(yCD\���6���*�{�|`$B������k��L.#Y��`:��δ�,gu.�W��9Q`��`��Q�?��~���{�������[;��*G:D�_��Xw4M ����tZ���P�13ƛ��S�m���5��jAA���HM�� ,��\�Fr�s8�ת�~���o�]qy��Y�2	�I?̃N��>�J'���[��p� �g��'����	 �9y�[�\�U��,$
9[��:{�$=D��I �t�;��ꨍ�]9s.����΋���Z������&���:��GJx��`����T���muT��Z:��N.U?�
O��b!6w�'�������+�lz|�[H>�Yr�̔����7���?;�e���,zy�!Z��X�<'~Mb'�X�A���u��e�)X���x�A����r\�Y�b}��E���%���*Č�cp��\ܥ�n����O�@�3촇I��Yu��;!��W ��t�c��~o#krź�2�4���C�.�l������O��7�sH�ݛ�d�?>�=�SG�D�7�����$��睿���]��.�bx��-�>�EZ$��i*u�Q���D�*o���]����i��O�2�!؀#)���T��K�6SM��^}��DҾ��uIF���"- ��L���y���K(��1�'�.����`��Tc�׹d�K\�]�w�SR5M���rW����F�u^��ߎ6p���7z� {��MO�	lC"���|Α�bE۠a搿��""�S|��+ݿ
P�G��VJ�aj�M�w�����c`�)�R�<�7�C�˛*�Zu��.�e����R�{~y�{S��2�C��-��p*��P^���?��h�1qPf�uz�O��٢�M9�
3�K�O���J��b�I�Y@�c��+?uK_�yˬ����N?aD�3~���R���t�Ʃ��t��1�q	Q��
�=}���럊˵y��h��|g�u���g�Ȯd���q	ڟ���к/��θ6>b���Q ��,�f�]��ї�E�m��|�mޛj=�y�D����<���"��%Z_�1S�	����7sA���؛����6b� '#�Y��˻ vTG�z�	�i���O��R�.l�f�t�F����HCҽ �A`䳿p����`�.Cȗ��zhJY�%_3�2���[AR+�����ӭ��)���ރ��0b��yh}o�Y��mx�LH��s�}�q7�ϧ��ls�=٣%�ʁe���ܨsm×����T�%��j���S�o�.>�'�u60<G�j��Y�m��+�Q��ɦ����nD��co]���ʓ`��
i��ޥm�@���@O���5U*�G|O黼RK�g��t>`�Oŋ�%�ZO�!{I'M�݊�ұ�PWV�@;������� /���/g�Y�U�I����1�!Dw��l �G#ЭYu��¶r�}a���@�{C�ހ���iA��|#C��?j��?�_,M���"�z���񭧘j?���e�6�{�=K쓖-2d��m�� �y��po����(���)l�x�,�x��ָ�1!̞�¢�7�/<�ST��6R�U^����rQ����/+V#(^X�"��E�ϒ*F胼�0�2ߊ7��;����ƺ��Iu�NF@ԣj����r�B�bC�2h<;C���"����ڏPds�Yٱ�W|�c�,��+�g<��������9u�N�'��[˱k�im�� �vq6Wg�_�$���h����I���.Z��{�lL�^GxK9�Z|�=��Q��/��!���/�-:+lm~�a�4l�+xƆ��i�T�����ѽ�7���(x�8�1xhU��&f�DC?�^�� �w��*���-p�������CX�����_�:qn���w��_k���u_9Qe%v�'�cf�b���F�u���G���-�������~�?ֲ�T��P�#sV��Z��6���=��r/4K:���0+{4ř ��\#��W��~��%3���[�R�6#�٦��:�tE_�_Ͳ��g���9x�;~á�>�ƁrRAp)��LC_�6��}��^k�����'(1Ѵ�!��&̊��S��<��j3�G��@������a�#�sjқ��SϻI5���aQG[�{A�5<L���hLw�-�'4���b�#$�/J�6���s�?��	M��xH����"��'5ď��P�j2.�9b��{�OdL`m��Zy\}��@¤��a�(f��?>DTF�E�M"��'"蹦�1�r���a���{!U�Oa4	���jO��"m�Q+P��Qṟ�sߩr�à����_
��P�?ss��4�-7���0��@�ٿ��Ɏ����EOp9"}�_9>dY*烃�_�4�h��4OH ����تd�na�X�K4���HݫoN���o�I� ��[�kh�[̴FC�o��QQR�y	Tvj���Z���CE}О�]��Wo5s�&G��������!�27��3��Q^�g�[�r�mHt48�S�f�.�P=��-�xh,|�^���6b�MGu����F�K� �F���HՆ�;>&o�3�)�h3O�0�3�;Yϼ���VZI$�0*�����x���k��'�)����O�E;�������F�jc���0�T��4�@9M$x��!���*� ��A'-D�x�i-��nL����p�X�VfI��ZAc%���J�l3�J5�b]�YݠȔ�z/��(=������q9FF��\ʥ�����*|*m=\�j�Ů�q|w����z%tV���}��A�a(���p�@�,�Y���i�VsR�Jcq��� �!��Ż�I5ڥ��0.�����)ʞ���h;�En�e\t>�͎� �(|~�`ґ�|�n�1eΤ��NݥHn�l���0�2n%�Ri�s�H���ښF���+D�\��پd��z��C�Q����=MsZ6<D܏�t>lϿ��6i�I�w��ST�o"�4� �W��R�iLuMD뒹�A�ʁ�-��3�lM�t�\���1���|�����k�>��ߥM�-i\m�o}#,�_�{٨�c��0��|C���i�#�1�G4��G�LE������qĊ��KǑ�,�D'�h��$1����KP ���o<}�0������=�+�P���젡�`d��>�Y��<��˖����Qܖ�O>۹(�����:�w��u��i}�ۘQ�jIn�B�p�^�F�\�t^��i�)|�[ކ����(kЋ�mF�@�k	���� �<��OBh5Ԩ<B���?
�G�A�����1��
vib|�-S�n#�E|��c���[&��5Wp i��Ӑ.{��r�h�}���`����	���Y��Z�)W��>#����E���X�f]$b??����I�)T�+���q�	����3l�[�-8\�t[丩��Y/�PS({���P����#Q��rwy[�Å��t4��@%�Ҍk�Ŋ>��
�_@��*1�@��-wi-d��4JJ�nI��;Uu4�Ʃ���
H��L�C1����Xh�tn={�b�w�!'��MM���=y�L��#�T�A����G���+�P������Fj�N�>@�]��&���Q�߱�KJ�m}�q|B�ߴ;����\A�`*�8 O\|��&L{��h��Uv[����
�L�]t���V�������4�_>���e��Em5z�ǞOӧ���-�
l�#ᚵVi�H��4���9�%`R�� H��o�����qB� Wz�_��O�)EaUv��
����*�4�M|1�yZ�E����;cx��srr��>L�J&��L��[1�mf�k�l/5�K��z�đ���b6~@��eԴc_�"�:Gkh�b��'�[$E/��P��6��U���N"�Ұ[a�x�/��[6��EK�eW�[�3�!r�#���jj ���Mv��&1ëoL��~��kt����i�ޗB�7��8wA��)��\�.��cbf���q�{�>²
�:�F[Z@�#���Wmh��kz.3�7U��� W��6T�1���ЗxI�!���&�����G�R��#���>��^�)�ʽ$~��$2q��_oy|�aot�6iڠDj��枏?]�L�ds��Fz�J��^zQX��ۨ�A�t�:@�@6]��&��S5�<`2j\b36#4�;��K�����q��`0�j]�c��3�|����i� �M�����J2l\�*ix���?1d�O�������N�p1��G6u��ob�);���4^k�ȡs0����%*âZ�=��=�2����t�=�F̽��� PF�T?c�ޟ����!�un�-T�0��כ�`����J��W�Iw)��%.R� ��ڇ��� :� zP�2�)$*���RY����[%A3 `�Qtp��DYQl��i���Q����p2F��n��P��S ���n��z�.-��ߤk"��$Ǽ���UBQ,�*�d+����E����vm*�K/;L��Rls#�Hx���j����/cl;��O�i�"-�-0cAS�X�}���"؅�����`�S�JǺ�zH����.L��s�r�j�!Z)�V�fzs��e%f����5���
��+#��6�{��\q���`��3iF�lb���3o[�:Zէ='�������􉙤�xd
^;ؑ��]�R!ŠY
�Sx
B�=b�5��u/eR`���[�l�:+�O	�YG����:s��m�o[��1�5��
�D��2>r�x�����kb��KG+0@�P�pb���N����}�8�-��>!�����6�^�]e�$��<P��c�0��A��̙�
he�M�`�]q)55.#e����ƻ�o^�3Y�!���VD�nAU$�546"�S�۳�MpЯfF!��������C�����15/�"S8�eiOC1l>���rOl��Vi��R\ܤ1=���]�{�T�����ƇF��7�re��n!0��=��n�pO-t;�'�?oӉJD����
]�J4��K^�_|��q�	A�k[��V��r��e]g�\�[�d��{���x�!l�ln�:�\u�;��"xs@/1���MQ��(KT|ރ:#�ڟh�<�R1�X�<�0�B���Gf���=�`��a{>�Uz�{s�b*��\�V�����ߌU��C�(�+�������u��7�ݗ�u��g��^��
��s��!wO�l��1��9�	s���.���V��sD#�+�!�n�k��;|��7�(P��"a��9<���8�&�����=^���=b���q�S��� �	`��\�5�3�R��=���Lע����ݯw�k9]'�OYp�C��}�o|���/4���]z�����M�m�V^�������V��bu-����2�2�c����.2X�<Z��w��4P�4�jk!���$�2K^Ŗwn��b!��{�����%�{.�E�ϥ�槭���HWo��=��D�M ���W#�~T@o(�N�I������=�P=�hl���9�Ӊ�/�,�� F�5�XO�åZm�4+���&sp���9.�LǬ#l�� 78Z旙X�N�hyw��A�I�{sؿtn���`�˻��xo˔����l��g�q���}��L��J��M:��]��W���U�&3�M��hgf�뀕�so����`W2���V%H���|t�M����]w�O�{���O���6{@���nt���<=����5���p��"̠K�WrCD��}�⊧�¸��������z���{+!U�nT{����m�6�o�w���ߛ<�������8hY.�Oɼa���i��{8r|�AVS�y���!�br)1�&����X�u8��jR�?`*t��R^	cϋck1V���o�q�ĝ�,ϒl������
w��DJ Bh��=s	��nn�y����v��z�b ���lp0M<֪��\�j"��KnkW�5��IDW�=�7��i���$�ԤZ��v~/�v+���(Ȭo��w���;}-� xT�>Y@՞�(=3k�m���R��S_?i��D�d��R=Oh�h�ʘ�ǖ6u$PtK9[�b&���c
���f�p�yma[���U��\��1���,"�G��6_�̽H,�3�u�Li�� _rsG��Vo�eaS�<��0u����,�����3�4���y��/D�Ǒ�Tr'�����n7Y�'5��LG�4��0O@���P���WIۘ����"��A�w�&�3���O Ҁ�<%�:�,���U��������>1$�`-s�t:�e�.��/i8�>Vߊ�幂8�O�qr��,M��/�!wrs2�cl�	�r��e9vu%�ߨ�J?^0��5�`��T���Rϩ���:	4Ԙ�QA�-���i��BY��]
��@�&I��K�MxO!�z�`�~��F��،#DHU�˽�B��h��Oӯ�� �T`��+�ֱ��Q�w?)���g�R�o�q�ۊ
�8�r���`4��{�I,���L<�`�N1梿�ݰg3�4|Ϧ��9�ɻQr�d��x�VP���~�K{c���煡e,��P�v$L�u-t�*w����R4O�s����u �� {E��v½Gb@�˯��Y�΄r�5ÃO�m�Nټ�p�u�b�Y6d�s�kml���t޶�f�(��j�(�؅��Ȣp�_�j��8}`�>���������l^ʆ�cS�4��%g�ܿD����ߦ�f��/����dĹ���ۻ)��Ǽ[o1?2)���e����]�yA���ے����ž��x��MZ��n���{A���Җw�P������tl�S���m�1bo6ᴓ�WX�L�"3w5�~��Ud�}�<y��%�0�OX'�����
��\(��z�S��,:�&�&����j�,�&u��>&��NN�G�!��_� I$�!8;A���,��+~xk>N�0�O��f�����@����IGm^��t�D�S�����8��]n�&#����f�n*��D�@&�>�É�f�l�ʉ.�hׁ�l����c��	�c��ϙ`�C��%�����i�_��� !q����˅V2ÇhD�jD���S�<b�xGcH�:X���q�aI��XZ9lA9`ئ�^����K70�A�\B;�Z�9�!�|CU��Ɵ�9n�i�5�QeY���䨶 z#��ڙ�>���!��k"����SQr��K���w>|J�e5�4��*�k�J���'��*���Z#�}��nj�J��L+��w��Ā��隥2��M��TR-%�D�b����7��Rv^��DV����hUw�df'#�+%��yu��ȍg��q�I:0E�F��"��ɍ'K�f��'ʹ���!W,YtB�LS��	�E�@F�e�x�hPgup�;w�YA�y氈e��p�f
JGg����ECC%��	SJ;�,�2�}������������7�o�I�%������F�@�ᵙ| ���ީ���v5�^5�]N=�qji�#����OY�t��r«����_���P�����%S$
�Tz�1E�Y@���f���1�lS,�����n�0�]MP�s�h� �&�D}�y�^�ۋ�Z(�,8ߋ\[{��Aօ���u	�%��J;�W<��*'�A�-�m[��ץ�m���kۃ)p�����I�f?ޡG<A�z�	M���jM��k�`O�SV��CKT��Ɗ���\���T�)����ѱ[f�W��?�޹%�O����o�r�����
�jب0�%Q�n>\�����gc�7�Y�|�A�\
T�י �o�$��du�KS	��6[�9W-��`��f����{��Z��rB���I�G��z;,�U�㳎G��9-xɌ�\<��7����=�����>ގ��&�+`���gj�-������J='�n�'�ɤ �<5?J�$A� H��k��~'YZ�D�{I�~Z���*���̊�d���ܴ�f
H�����'1�E��h1���k�qc�6	��+q<��!R���Cue��
͜���V+
;��Ye�¡hV��B��|� �t����Ĉ�i��0�����	՞��߹q�-�����?�>��8��g���
6������N��0��D��}�@`�@��=.0�Kޠ���6��+h�|�C5*��HO���ۦ�c�05>��������i�^!�9 ٹ�z_� �Is0+�ep�1S~Ijݜ�	a,�Z������Q��(���]�H�����ʜ���7�����2e/IE��:�x�ȵ��F�[�ђ�}'������0p�����������2�/��9x��kp�G5ʔ.�h��|-栆M
���'�9Q���E=��$;
-�ާ��n��A���f���&�_�[%��l�[O�$Ҕ;I�_�c����u�Ps��]2�C��N���g��]Ik|����8@r���	@P�.�� 3P�V��a����޵5��Hf"�bc��I2�����b�@!�D�g<pd�
gxK�y�j��� Č&GANj�@Vn�r^+�~�%�ȴ�tA�'�2IMH�z��F<0���*�R���^�z4��.�6�:*��Ժ�)OAl���Z�]"(�����؀�Cc)�C�~`B�sf4ͪq1�"��&��oL8�vV������I�{X�������yh�[ �2k�~�k�J|�I�$��q(a]�*7ͫWb�����&��.+��cq��~ҊŃ�ª��
��Ĵ?ה��=�kd���*qQ]ꊳ���̡|[�L�����T���㖯i	����� 
�����iH y.��B<Ȫ@�nJ��c�o�~�l�����@�6 XI�e|JI!�<�Ϯ�������縶9֪a�"���E�˂^ ���5BfwX����`A�	���et
�Ñ'��冢���Q�c�tjCYhY?��+<��y�)�a�� ���S�fE��[��m�c������st���ΐ�)�ʣ�m4�y���e��۳�~#!3�#����J�}Bj�j� �u�L�WJoo�P{�wM�4�BB�������A��A��[A��$E�h��{V������#=�/c]R\i	�S�,������Y�&SL�����������.H���4V�'}���Z�N�~Ź���|*3���q�����j�������SO�"���t��4�,0��bn�e��s��6�vd!l%a����'e���	�����=;Lu����I�DĤ�S3��=D��h�=t_���Q)U�	����	���'�k���c�Y�a�!	�.H��`�=�'NK���b����6_FC��Q�My����T3��T���f3�3��ݝF-���=/0ڬ;���Y�fٷ�:�V��RT7%���pz�~Q��/�3t���F5�nFX���Ҫ��z�F�/._����jNZ.�NGDi��3�Yw�}5qe!�2�����x�P�Sа�V([��Á�XV�"��J�M�R1R�Y�*^��ٹ��q�#�]�V6XB�[}b��~խ�[DX��nK��*�a>B2�e�ž���7
dP�<�ؾ r����~j\��=��fC�wQt�E��򯪡���ax� ��ԚC���	<&��+0��ۙ���Og�����|�k��8ܾ�t�;����¿�r�(��@���r�8��_/лHؕg�%)r������!U}��`�/Fk�S�S j��D�*ϫ��p"�Ak>X��7�#$\F�ɍ�Ξh��,�k�kn�78?{fc)zn����]w_�hf�T�=�O��1T�&�ͧ�`��룆��QOF��p�qL'���?e��8��G����9��/���h(��_טL�3�J�j�~�RS}��$��>]ɮ�L�L���dt����h��S��bu��h��[�#�Q<��}�ZL������ >���<�g'bLkJ)GXbB�z���^Q�yw�Z�*#�R�k�X,��������Ƀ�\''IS"�q�<H��4�a�=(����J������%4�Fb����U�r����k|&8Ɠ<~�U����H�8��ie����ԥc̉/���b����!��4':�y�9�E5L��uh\A��1QQ.�ϲ~�E��L�/�2?���M�|7x.�D��0�lV�؄�q����U��ԨD�*��+xgϽ�R�}�����6�X����<��2-.�� ��\�%w������|	%��|�/���^t)� �x���v�zR�978:,};>��TU+����[��(Tf6U�=��_���`����9���G�]�����t��(���D\�3�u�EmjZOm��Ĉ��3�ʄ]�1,U]j�p��_V���P'�)3^K��1^�0�M��c0sL�:���;��7����`a5�䀯��6@����S���P7�#��mZ�!�Ōx 2����a|�؇�@�@����v$������$�;^�.~n[I2��92ޕ���H�+��cI�dM6e��ù3Ut�͏�G�g7���!�m��z�s�~��-��L~��@W�֔�2g�ĕ�)�K^�Y��4>%���<T�jdd�F�:�k�/��t���9bM󑞶��:�/O��t�\E�0GP�8�J�:�0&�,��]����g���_���6���[�~�oϙ}�����0k��	Z\�1���Y�UES_��%��A���M
4\S���Ctl��"	b��rR>e��7�"���{���x�fm��#��$��Yt?1�c��ۛ2B~1�l�q[%)�Ͱ�y�ky��fz����X�u�0�c^��23x;����Άk��%�K\���f�G;q��M*F�m�g7���xdqz:kײ#ot�B[��P����# S�I�� �4o�6�:�I�e�lu�-b��`�!W����W����^K��:�q��\��~���nS,��� @X�Zo��U7��qL�mmC)3�8�m0cHͻ�Z�O�6��ݳ��(�!r����q}_�k���x�G�׫����ƒ�C4��'!&����%nl��]'1�^�U��1���R*� �;��U:0&0�$�M�0|J���ao�AEN0+��X���J��:��F��}�2�]m�t���9��IH���L�d|�,?cS�qv�Ո��u��y�V=[�r�V�Iw=p��b7��mKk�y�p��������9���*��~�B�<N;JQz�;t�)���L	lćf�W��s���h���3ϋ7ISh����2Ւ-чQ�w��CN��~ �:b+Oͳ��QT��5�*e#{�����rq�v�Z�Q�$�5�H��^������P$�=�"��b�)���;LW��/̦�x����V�� � ��j<ՠO�&s���[��G�q���q^[/b�Wn�ӧH�&x���?5wie��l���n�<�m��R}F�/h
��r��Dh >��������$JwxM
���˿�E���=���y��OG���([kr��U�>�UI�~;�_���'+|# U�#��ɉ:ݫ�Yp��� -�_��yX�[V
~U��G��\����#����9�G:VO�+| Xe?Z�U�6�k��=��Ǚ>4	*�{�A-��#�ԫH�bjp2�ub墀��ڄ�y"��5��v)"V7�`qĳ�N3@�޿+u�oY ��>3B��@|����dp�����n.u,.)mq���P\:����0���;��/���S���u]��O�g)e՛�����M��72�>$��47M�o{Qg���m:�3<8R���Y?�t
����$���-,��X�u�/I�=����`���􈰁�y/�j0w��4*�U�{"���!�
�x�2$˸PT�m�௤f?�>k��!�'�Ka��k��=��v�я	c�Zú|X���Ku2������ʭ���)���������g����'(ByKwY1.۰�$Ij���!kToMc�O ,~2%(�B_a6(5��E���� ��Kw(K()}\�ŚE06	ޅ�N?���g�����@� g��ͩ�c�f���� �M 4A��H��ŠY�F~_���#p������B�#-+^��3E5v�Q�Z�є:�!�.�����r�~���z9amzn����g���u�k*1��8����7IӪbp�Aq6����t��ݚ@^.��8�G�H�p�b�.��E��]����4W�^�^��AZ�Gx��6��h����r��Z��#��Y4묀���U��j0��"E�L*v~����B�)��>ь�Hg��G%�`��.�$u�����i�ú�		?NY�zr$��'��K�H��4�1ڪ��S�q� ��+�h%+;�m�$&1`2��_���g.-^݊e�bSf�B:z��Րjz��
;&����W\��' ME!W�^?䇆�lwo_��{D�~*�c�=uq^�����>��c_�s+��XƜTj�ZmX`���4諤��	��{�cS��͡�6�Fk4`��ʖ���1���L� ۭ��*�h�^�m�^GEK{����s��ȻRѧ�����k�Ne�8xS��nT%����l oE�����/�6�I����@G|��k��T'ov�R�~�Q�	��Q�$&��_�X�R9�(�\1V�u�H�L���ӠD�*w�����p�/�i�)��5Sbv��$	��wLR0(��g�w�
Na���Ƈ�����	�Az�=)3��8�R�c������y�8m	{���_�_t�<�'Q5�ej����:����/����&��T��(�!7�A�����d�yH]Ev\#���?@�<W���J����^q��hD�R˫�UL����O:�\�U��<������M�2�@5mD{�]�_����_`P��B\���?$v�=�u�n�(#x�P�=c;�l�^(���!�6.�?��U!�s�ul�c�W%Ÿ�6���7�;�5T����eB�ܐЏ�$su�5�b�Kr��q�Qִ[�@����4�4����s����fҐq��0%�L���ڲf�x��rS�.�ˮ�d���6@���3����6�Դ��@��w���j��E��D�R���G	��m[r��cr(U �����s�+oq���cϻ�<>����Z�g������
�itY4Ty��Ҟ�IZ)�ws'�̿\;�X��qdWR%����Q���m�Z�ַ=i�fv���J%�|#� ך���"�G��%W���k����%Χp�)ۡGC1�ǋD��,h�	J�G���^���� �d��^���_x�Ek}�����*ug��H��,$1��O�$	ov��:��g,C��9��%�2�#څ��R�Y����^�:�| �UN&��t�_g�?� /֧�	d��F��.��)���x1��[v�|��d�P���<�O[T"R7K;�8�x
��˗V|�hC����������*�~�~ކf��R����M��b	d]��
6����En�ٸWÛ�ȳۭo�2�� b���Gg��t�)�*u<��
+���+ݗV����	n/zt��c���i��Wi���\�@��d���(m�F�l��F\�3��@Q�P--�j��z��72�N�5���,�*}���(�������)t�&ͩ�&�~��v
�ĭL��d��`0�����4<;p4�w1=���N;O�j���m&g���4~.u�GT�S��	�e~<*�NН���k4f�Ͼ�� �d8VWA���ME�I�WD�L:i���	�xwe�q\�ߕ������=0衫��(XA�6��+�v~���&����R�,�V $��>�TQ:��e<>a�-����<[&8O�T�E
¼b�z��eX�~	��ޥڿU͉�6�P54�],�,Q���Z�����'�G���Hx���6ê.-d4�1�)b�~[�o�r��	;�&��ã�����t�\��B����f��ݿl&�X� ����b��p�wO�;�B7I�d�GQyVL��l+g@�tHg�忂Luz�&�	KoEΩ���@g�^fU��;r%�������ȿZ@��g�,7���^�IM#H,�J�R-�IY�`���9�/���ݤ���s�~C��V0c^��F��Pt��v��m�4���z�VY�rk�qƉ�@ �ۿW�y\�o�<�r�m�#N'����~F�!��È_�{� 0hb\U�����r_�˦~��K�������a�z�k�����R6"6���q��N4��Y�a�������,��НB��|H�f�V(����c�	�B��v�6>oی2�!���Ax�� @ޚ�b���k��E��9t�Sѝ�u����U�7�n�/�6	�����w�y~�_1�X�����p��\��~�
�d~�t�K�x�w�M=��r��.6���$�B���Wb���z� ��-0`�[T:��:�_{d7��?���M� w�c��t  ���I�"a��H��k��wV���NZ�I
 �/��pផt��@�8��Cmr8#�ipԤƩ�����4���~uGC��n���j�\#S2Ѧ�I@Խ�PT%|�Ү��
���sͷM����,3��Q	��:^$bK���Q���+ZJ�Z�+k�˙�,�y����E����4�0D߄���!���j�{	ME��T2�1���P���-P'��D{=�0Mr`Ro�������F��ڶ��
��}���8�^J�e-��;��} B=�3α(E�˃I<ih�4tӁ�Q��ΡS���ݥ&n���d�Y�̏��cO��.��`�=\�N�&�IUj�L��ݶj"ưL���Z�+%��΃���;!����?))�ΐ��q�s��-^Xks��}yQ�,��t,	(�R���tz:����\�ę��s��3">��:�
�ji��(k~�d9��C�����C� '�)Yk�w���6�ڌ�l..߄u|8v�[�_q����>Μc���
�L�LB���kOiN]�܎UC�}��#&H��@���NI�U��EX�e|��2b?�dҔ�W^*]h�G�������iG�M��%���x�

���A}�F�F�m����4��6���^Iy֣�δ�!��;6�b���o��Y����F|���u�r��N�x��`�K�s}�ÆH�'06x������#@Sב�>(]jM�'�{3v�l �lH�6��o[O��r����d��>�"�a�"��I�r����Q�Sa��t���v.���pZ���_Wf#|�1Xy�
�C�Sa	 -$���q`_�Z��ta�˘a�g�4�939�[���09^��{a�;Q�ؤ�R�S:��ry�&�Ӝ1)r��T��r"���%�9)��ڦ��%p�J`DZ	���p�6-����l��i����1KJ��Ϲ���`����Ӵ����e9��d�|�Tх���v���"~��?-�q�7�L��۩	����^����C�M,E���z�����#��A��E��dV]ўLc�=/a�XĪ�K(v�#�t"���E�\o�#]��M�����C�,A>z�I�으�Q�,���rz�\�}�D��<���y�!�R�R�+��aR1VQ�]�!ʜǨ�?pS�zzׇ8�P�M�����Q���j�'��\N��fF��U�2B�]Ԥd��<�������8戋����Ә�<�j?Ry�͂�7V��gs��М$����o%?tҒG�ҒN��3�F
���pE'JA��z����bk��5:�\���:�W:9+l�NJP�َ�-Co@'�'��͌���4пt�����GJ�_ޮL�8Ĥ)j0�G
���{1��w�9v�$����1��o�����{�6�0�\,�<Ui�@O����-ߍJ󏀭�	�o�G�*��~��Q��SXBQ�+S����J�rW~�Z�6��q��Zw�ۅ��'���e���q������;��!=���]H����g�<-��?�`q�4�[��u�I�OǓn�ːЮ��������{���btB&�Z�����W�G�Kɡa��<�ڕ���#S�}��5Cl{m�x�'^ߎ9�q,0)���e�u@��_ٰ��0'~j�5#6jRY�vim�.�D&ѻ�ƴ�@�	�)x��'��g��0w�6�W٨Ey�3�Sr�^U�5�KI|�eD���N�t���+<p<��������C.�?�o��D�6IO���'�*� �肮�L'ܴ��ez���|��a_䍰G��~���2�,x�3��%ړI0I�egs�"N �����,�4��`�����HrE��������!�bCgV����Ǭ���E��ӛ��wʹ�˔
6���y����K���~���
��tLp%��.�Ń]c�L����$��{��l��߻�M�,%�z=1<!(�Ü㑲�M���hz�6������4�-]~�Z!\�0�
󁭠m�nj���=�-���M؍�R�f�xJ�s��]�lmhǛ>���gd��X�F�V��<��ZA��k�WW�7=r(]�6�K���3�Z@������o��xgPP|m�E!��0�	Y_�p�]�5�8�Nr�����J�k���Y ���4��{����]�6L���LT�S[�$�V&�w��{!ET��r���7re5b��3ҼzU0S��Ȥ*@�b���Y{	��} 	���/���C���
�iL����5�EosZ(�ؿ��W;&���q�v�ë��:Vv�C��A�y�[~'���h�i�(zm��Ρ�}7�э��1���|�3��-�턁��4Tço=�8VL�{O5��8Z@vy�q3��Y{��x�Eۦ�DƙN�:舞��0����z�$�-��?�?゚i�?;������G���s�e�f�dH�ۇ��UΪu�"h�g\���,Y�N��\ vI���b%Ny���(Xa��R5���4�]ܣ�H�K���h
2s�S��摔��E�㬎�=B=jlϾ�|�p^�Aq�}�W֌��Æ�UG*(RR=6y_�b�P)@��#d�_��)q��$l�:Y{:�;����� 2l�=?��iF��N�ؘ/�ɱ�9�����ˁ�Vտ�"턣����vgu���ơ�&T���j?9u�򼠈/���S��W��8�O���R�h(OTU)@��DE�x �\G!Ð���h��zX��?6S�!�DX�
?95!T�Y�H%��(�
v�A����ŧi��
Q�v�9��Ej0/<�@�D���j#�8�� \ߔеx"�1���C4fZM�Hv�P���k��
9����=(�t�aQ��Bl}�%�}��tm��Q�:� {�B�M9�2�]���`]�Q�0�����,zp�B�����h�M!V�^�\�p��L��JC�S��DUJb�g���Q_�Gr�Rֈ�(ߥ�U�,��s ~��V+5����߿#�����a���h�W�*�O��Vz�{��UZ۳���������#�����
ȸ�Za2�S��VF�H�ͩ��m�"��P
o�T�O����ٲ��*�6_�Nni���z$	U���sF�����>[���(��O�!|�����e}���:�U����������dg[Z[�i����2�w6S�:�D!+����q*=�s�b������W�g
��9�J���[�U6���[0�?��33,M.W6��ܾ����eEEF��Q����o�䳟������{��cu�G�v��_�N���̱O���C�5���)�C�|"���'U-u.yQ��wn�uU<O
�Ơ6o~V[�0HJ&�`0.?0!��
�A�#�ɮނ䞪����\��%��BA&����!w���ԓAm�Q�z��XJ��u���ɳ��9�x��]�,5�4���&e|v��ׂ>U����mP��Cwֲ�~TB��k��$`����0�t7���T���2�,a'!(��_�S��C�;[���A+"�s#�E�<��X^��=��G�;gz�����sur�վʾ��Iۄ�]r�{��R~҂+������v)�x=;Њ9�s�t�b���_��ɡ��X�@߄���P�_�D#�E��
� �z�������5l	��\u��7-�ܦ�C���8��e�� �hͭkH(��\��2�_�o@x����j����Ӂ����{����'{x(	s	��T�����Y��H�5����B˞�ո��z����ӎF�G!�qj�F��ܯS��03j�v�D�@�������؂��p_.9��.�O�mj8��w(�̈9H�;�QU���u���4��;L�;nQ�e�"j�����Z�SM4��ntL�샨�O��ʊ�DdJv��]��a!q��o�E�͖a0%;^`�?��E%� ��Ƌ�*��dhE��.�{�)4���ܷ�'g[�_0΍��t��GpR�*�ց��Sx��a��Sx<K�s~('��!e�5o̖:u�|�g,���fo���X#����UeN�"�`��O�J+��wŶ=5�Ɍ��f�Gi��qb,Xi���e� �Nt���7�%�F�&[�'������:��S�%T�<;�g��p���^5⨊�{y�M��փ@�Ã�oJQ�,h���,� G�Ճ��],�,tg����t�]5����ns`���"R˽��������?O[/c<�j�?�@�������l\����c�g΁Ћ��qw
n'pɺ)QF�G�B����כ�!��sx�>^�zb	4M4�Sj��T���Z'�1�m-F�r�eږ�x����)���W���W����j���^ϒK����ڪ)�C5��7	��w]�rK�6�" �v􇃂W�<�������\� ��l��<6�$d�+��Jk.�O��B"����r����P{-Bd��2&I*O�z�m�&"c�zD	��bm�τn6b��A�:�i�d[�H�T<�j\�-��U~��V�;��4������)4��N�U"�I��]0���+.�s�\���jY9V�V*޼$��@�>��X�rr'���#"�E�K��{u�ND���jҸF͈"�v#s��	K��&p��'m@?l~��Q~$���=�Y��M�Ԓ/
�_�a���}Q���?\���L��/=��(B���W=.�"q�q�F_���Ŧ$�q��d�����+�дC\"{,N��)�7q���'���z��j}��X=�{��H-�'�`&R1��j�C�H�6�@Ího!�r0my/����?18���W�a���w1���wo��݁D
o���lF��e}v���3�5f�1YD�k<N1�??����!ݮigl�3l��"﷬FD�}���F����m.q�B�M+��Sv
"ؕ�N&p�:��dN˘�~��\u�L�q8���	��CF��gR�
�n`���&��_yha��P�*A�Y�˅��Xt���n�q�q~?#�e�}���9�r��m$s֕���5�e(峡�ɓ�X�s��)k� p��ed�J>x�Nt\�-�*~Gѩʾ%R��w_�M9�9i#{{��Z�on���B�3&
o��@�5��<&��6�fw,�LF���nOn�1�ȋu�؋e�4`�*�v\�~��x|��N�IK�6�PҐ��4ܐ���Wȥ�L���9��ͫ�n��>!��m���a�}�w���٢�̢Wy��CX��0� ӹ��0\�E��f����!�TOp�g�{C1G�-� �_a��J=�/`T������_>�Aj��4�#�X���Q�&���G��ߔujުcY�����?J�m����G|�C �k�m\��cBn���Zy��4��]�Jȵ�/��IE�����������������b�!7{4ɏ��Q���!��D�Hi��S\L�0���Qf^�~s> Ì���6a	���[@�8�=��/��/tտ�����B.�>�&�� �T�*�>�������~.�)
v4'\�{����^N ��5����E�E�q�z���Sq���czW//TA��$���"������gõ���oɹ��'����M��/%l��f���桒3u-t�d/��se�������e����_�T�zɿ�1�JjѲ��O�D���;GԔ��*��EģSX{��1��UL��ę�WG|�sx���<ym,?�jd���Nqjd]��R�*�;2���Z��L�;�7긷f"��[*`��cE4�A�
�pqJ|����V{�p*��V<v���, ���H�-���;�Ҕ�)RR�s�������xp�*�wXn�Z�%�Y���A_-�����F�˫���b��z���B�!�U��l��=���bK"[���E��5�\��j�_ѣ֮r~-�a�5]����.ޘ���鏱:����-C��v#���	@!�o��5�B֞����<��&K]�<�,�qi.*��B����eo���h�0�]^�:v{�|����Z�Ǣ-W��q5@tk|����GT8ՖB�!���ȵ��B%���M}��.�ߌ=��MVe��:N�;e�Ҹ��h59�c�( �����|>����)/<WDl(��7ҙF�*�/�����J����������'��W� ?�3�G�aha�I9�sm7����E��?���8zȁ�����LB�~��&/
����Km��h���a|��UB��� �I��g���0N��-y�������\�(C谙鐡���4�{�y�jC��6ބ��/��rp�PkE1}6[�Ց��ܤ�=	g�!�a�,�e�ʽ�4���&�������NHuz-�r�vJ�1G���b�^9�� TY��C��F�	H�0�I�YB�R'
��_Ø��c��9j�ۙeL �W �fM�$��Մ��$�xgջ�D((-�#�Dl�+�������ԫ�4ת�>�@xx���Fju��G��)�D���!���m�sRv�=�4Dl��谜Lo#���'��  ]E�q���/���\T)I��"���ט&�(���m�����=�^)�@ b�����xZ��F�_��4�B�mL��lP�ߞ{"E�Gj��I3�Oj	��<�܆|��ᄩF�y��&O���`
j���>+|��j}qpAf\=��`���c�j=�	�>�,�zK�A��>9�59	A���6��v����a��R.~�XӲ��t,�sx�]��*[qN�bk�Q-R�/+~&C�q���v�����F�Ч6?�e}���.) U���c�s��s���{�a�� џ�r��8{�$�У�m�.��6qO|��.��C�k�Zp�Sv�X[�hb�����.,����I�,��uE�霊�"�Af�xN�mX|X���X����Ig4W_���0҈Q1���+k�6�v����"]EvNe^o�d��2ߜ+󀮕Mx������8�;"�6ݝ���M�*���{�Jc�d���dL�TP�U�"j�Č�*�j���6��7�If�U�������t�{߲��Ќ��ɠ�O�a�;/!�7�#etU6o��{��Ua�<G��ד�{3	;(%��DxY������|N�:�^�g�S 5ϐ$ws�~���N���-	ލ��sUR��"�/��ܗ�}�\�mV�Z�H��ב/9�?J���G*�G����VY]���C�(��2a��ţT��f ue;���4q82��T�=����1���!�$m^O�ucF�u��o2G8��VgvEI�8y��S=�k�Ȁ-�xosN.Zg��/{�@����<q���&
������mZ�WϜs�ui��(�c���L>>Q`�`�z���ꇢ�ȯ,H�I���� U���wI��lno�%���Ò�����z�,�h�����i-�:on���8�s�'���~i��=��F�&��g����;�w�� �� [��R�v]��"�\���l�NN��� tWx� rO3��U�ܥu�OR@��a��mX)Ix�����W��ggt)d��vq<�7���.>9��������u�W�H����!a�f�Kr��� ��~�E5ʇ�=�U5�%Z�qϴ�6W�K��l�b��RS?Y>����s����$!fA� �
hMm,�^���~����U{ ��y��A5g�����o�J��(��J}�w: G`V��e�4g~���%_��x���DQ��#+�G.]bF%f�=mv(q�4>!W����ДVj)g 
w�܄jlC"�-9��U�vͰB������Ah��d��k�R!�J-����b~ki��ÎHS�i�a���'gXo�A�����e�.v�"�����D�x�����#k9�\�_�]�϶������T_�&�t��m	� �D�ղ"s��b���Ogy��Qn[��|KdC����݂��8j'`�|�X���W���̍`�w�BQZ��1��l���N̿�Y�f:�T�`���w�^+rI*Y�_�8��V3���Ŗ�"�-u:I���6s�u�EyFU,�g��k�����>�'/_�!�b��AޟTUY���`N��z����4���b�S�Ώ�,ҷ&4�%P5�$M`��(��T6�#�T�_��q�-m&�G���]�1nZ��>O��	^�W �W}�4�y+�����qh9נ�1��.*�b{u�U����	�s�W��\#����/���Yy)UA 3}ǀ��U�X|��ՒMMj}o�Sl�e��u��.�&��xX�QTb�p���(��թ�G���O�X��#�*�;c��f�͎gޤ��a"��8�#E4ldxxJ)��s>vɐ�͉X17GX�B����g.!�&���|��l���j�%N�x$٦��D6�(�4f,1�(�/�wB���I�Xd]P���Iօh����bɔ�ޚUoP��<	GV��~�&�>F�o_	�Y�� �#��>zj�ѻ�끈�f�Y�ٳ����4)�C�������/��;E,�fk�U �<ik	�Tl{~����NB|!s����3�Y~�d�Z�!�d��8�];�sY#�����[�F�"f��wI"L�:5�*�ω^������Mʀ8����y.]���D�U��D� ��������Tt����� 뾴����j;��p�Oud���'�b��g[~T�uW):\ �6�y��<����(+rX�<�]��"H�%, g�JF��rd�����9�eu�Ƀ�T���_��5hua�$}
?�;B�R+縻��s�]qן�60��sT��T ?�y[5�d��'����v���Mt%�<H�Um=H 4C�iid�C(��M
�A�|�4]Ԓ��E���Z�df�4�Y,��(J��NMKSSP���{�^���Ѹ�leA �*��0��Y�D> 6l�-
/��R�S(�H緟״��CmF^'�U���K6�jw4�52�r�g�׻;�yc���E�/�s�Ë� �}7%�݊.�\Ǵ�J�H�_���7��(���y�������x��+!x������z��MZ!XN�ND���dP�fRC���!�1Ơ�_;�>ġ<+d� T�VS�n'��|r8� �zI�3P�u*�+�C�l]����v�`��~bCX�*��<yL��-�W���G��.���Y�0A�I�)О�d�BV�@:]����-�Zr*���x4�k�{��#M@m[9�����d����#��F���?OE�Q�\���f� ��B�c\b+�]tG7�l�<(�!�B G�uN��{���7?w6QԘ�vo7������d��Wu�S��.#\(��Z
O� Y'��WY���,e�_.�� 0xG�Z=��_MTF��ۉ�nOYk�5��h�����my�ay@�:Ғ;M?w��z�G��rE	䆏�i����.�Áon�273�>��U����C���;M��Sz��oN�7؇D�z��1�����K�1�F��*A)�F�fE^�o�;�����[����k�l[Hv������I�7,�����n�����ׯ\��d�»�T�~K�Y�V�P!�*����2,��@j6��5�k����Z|E�5�?"Ek���6�����:aݧ�܌`t[�ۉ���e���1M8^�w���������5ݠlDW�DR
�C��+�E�����_��e��߄j�u��إ�)�WJG�}f�s� �����=ŜE�Mx��M1*ks7~�77�Ȫ� �!������x~$S�nq>?G��3�E-Cr�v�Y�p���>��Y*�=Y�Sy��<#nC��MaG.�W��;�#�-9�G�??��g��"N��3%�ʮ��W�I��_9(1��ߙ{�����;���O|\m�f�����k#���٬��/<Y�G\!�� ih8�3�S훸ĄYf�]5~�vm�T��A[kI:�������ܶ>�L���DE��x������tS�b#^_�iB�x�?P��ow��6}�2F�.��²#��r�v��Gre������w�V�E��'������'T�M-m7�9�o?['̳�o�c8d
�:�D�dq݃F��-�
��¹~��:w�T�sR���2�3�$.�����l( U������z�檧f:���d ��s}��n�*�z38��Hf���b��i��w�P[\%y)Ԙ��Y�ѹ���`x��=���Y�}Y[��s� �"&��G:��Y�^i~�WX��
�H^�5V��Q��h_�B���8j�9F�>���o'�X*�W>3_���2����8���q/�ȣe���ߔ^u�tͱ{hs�t�)�Qŗk��Q"�w�D���d��������=X�������t�W2�x�d��oTl����Y�H��٭9�Ftdv��jxϔ�1lq��\�@H�[E�̰s�'�G�r*8��wP�P�XjC1y*Sl��zL��@c�t�б<����uT�Uh�It������z/�ՠ���zN�`�`x�c�o�Zm'��{8-�c�d坑�,,�<��'v�����7�I�[T�|��X\"��*-�g�~���]�~�-�./��:|@7���	���������O���w�h�?C�cP�>�y��V����C� �z����_�D�*W�@�Wc�(���uo*B�p�����-�@��N�4.�����;&]�*�.~g��ź`C��H#3/�7m�ĺ� O�Ț����k�U��y�A^�h+�(�%IH�2�Vu��q�QB���hO9�c$��A��n�VT�Q�LzϭmP.R�G����qD�� �^��?�ͅ�q	lD��)٧��ch�!Ģ};���3G�9,��~�OM����H�K�l/��#�?C�n����2\�mn�1Q9��A�cn�_�PՓf��٥e�,��1��i���T-	�hh�窘5��dl���(���{��*�H]�(��Dl�QKV=kAM����i׾��T*㾿��K�#��|��D��[(U���y�,^�CsPӷbM���M������ݽ�����^x/�R��"33;��Er�>�vX�ӹ7�ڱ�����u�8�2	2x���� 
,C�@_Cˍ��a�!b��`���,��w�=���q�5�Do-�TfJ^%^i�C���mD$�y}D��N�\�>�Z��ƠO�b?��$HL|�(7�=�L�p�<_ŐJ)D����Z�I[���;w�,#b�F��<�{���Q��|�w)fa�@�N��,��e�&>��יR�D1ͩ] �5%��2��3�u�I�>
�?���S��8h� �k�E�@%?�1Ʉ���4;��P��/��a׷��+���������x�9}�TU��������N�j@!����{�[}t5��ԩ�ljZ���Ե� y��ն>�1����UʍQ�ˉKQU��%�jا\v�]��kx�[����
">�g8��D��.�\ �:U_+���tyЦØX��P��9�Az��[%�J�g�zq�!��'3b�ƪ�.#�F;!9�	�O�p�#�������#���� W�=�H��� �3O��z���J0�}��مx~:�K/����=qb�j ��U�T�û�F�cWnt*�[��x�������KS|�ݠ�}T�x����jX�T娞��i�v�iѹZw�^Y�9���t��ܱ@��>����|�w)��!$gk=
��}%�a�ś�ּ�{��ZMeH��H�*j0\��M�q�:�����<�GN��׹�bFq��5�D,��]g�>/C��E�������nµ�>.��#1x�>�#�&P|��2�8)��L�lUb�^'����uP�|n�- �n���]n>Z���k5�p����oQ�a�i�#��	�U���xf�w�aE�N녡�� ���i�eq���d)�^�-�~�;�È�F;p���߻,��l�")��u0㣭��j%p���0*�ס/#����l��uv�0�N��P��"H��<��F�[�8w_��yNe�ʦ��j}�c%x. ���%��E�\˦�	b����z3�9�.F��˨��X�mr3�k�Q�`�^�f�NBI�cs�^��Y��8��Kδ�\���G�'��ivH�@��̵x����:�u=K$�%.��$T����J>"1���m���H�a��m��K`�M�!"O����8ʡ͍��X�S4���R�;��Q�s�m7#�J����c%���ݟ�j�ǫ�\^kL9Q0l�R0e����n��N�� �F%	�a�a
����"C�Hԃ��(��*��Izxw^�e]����R�����3���/Q�5�lß+�E5�b\֍�����F"B�Y���V%���#�������9�0�v=���� _T�[C� ��>���JW�h�&�w��#\�
�˿���Q�Dur<ăe'MAp�����_�c�}-DU|+�������A��c�}c+B�d�Ue�]���ڕ�ˢv�_  �fx���Eo2�[�L�P�?}����j��8��?�/��O.�'9��٘���4���E��@�Fw#�L���	Y=��X����.��0K��F��se�GV�!�9�
f�Q<�K�zlkMƓ����ܴ�Yi:���l�Q�:�p��%,��!*e��@��OU3�F;M�/�ٝuT�eч�@�K*�4wl���_~�y	T�;ܹF/�����k�k��	�زuw
]�4��sh�$�˾M�]��Śk�)�i7ޖX�Q&԰�sCm\Ʋ`�\��\�Ҭ���9�Bnwᦇ�
���1����VJ�ȩ��Vb�n�P�2� qœJ��)�?��y������s�h	%0�؇�Vi1�J�����S��,���F�)"HD�s�v*���CsW�z�<��>R�����,a�/�ŦB�@�Av�_�=����mK
֋6b�@��;�����f��z�_���B��w�X<����І`A!��xG�����W�5���wSWr�ăT�R���Ӯ�RŒ��O�QW�#@�x���)�j9,}moW�����B\��<og(\���f�/���@�e�j�yB��)~�*��m�,��� S��p ޭ��
������L�X7��J��>l8>k�G>r��c���ruMJ��G j\/CJ��a�[����'�t�w��' 1�L��v��V������t-�&�K���L��{�ȉC���|6���}�;��h��|�w���!�7�|���i��=A�򐛖��4��~YW�FL�t�������x|�3=A�S|p/
�q2���6]�v/D�_��눠�=ܦђ
7��ń1Y�+�[gm;��a��R� &�L���W����� �K���ëW�ÿC�l��Yi�y�����JoBh�r	X)����Օ����O����<�݅|^w���G����e�^y}$��p�P��m��L���zB�z������r,C>�3f�g�鍊4����1إUr��V�mT��A��"9�wh��*E��z<�^�e����&��b�O޸k2�-�i���O���S��#������Gک�����;X� 4��nt��\~Q�g�E9��C��0�.��ES�������K�EA�֕������D-��Vgl�'�vJ?�����z2��h7H+��K�����K������:��}q;g*�GC��Q��)��.Ag+[	Z3it�*s����ڤ.����#��Ou$d/G��YV��iޗ�Fy�7���sk��O�{cu��n����xvcg9?��"��E�6�<	�����e9
�.z��#ff/ᴑrTD���`[
�%�ƭ�B�蓤��}WO�@�����d�Y� �&0@���z�Ý��I=��]�1�g//��h�1+@X��}B�I�?o_�z��|��2�4SPq�����Q�#>�7�H�	}*�i3\�^?���2���i�ڢ�����,�Ƀ����#�.ݭV|po��O@#h���Fv0ss�HN^��d%%�a0]�V��}�²J��e��Ӏ7n��|����9-cn�0����"~ܺ�|�HE�o���$p�d%�Uv|��x#e��v�J�:���_�;C�N�!E����9����V���3��N��y7t�v������gh&�@J�����Y�0�5�����5�A��#���P3�����2ۉU����Sm�@�I?�CJ$�*+���N�6~��af9�y����\��Y6�GW��+f|�q��k�W\�?��`'���af⏀���RwP&e�(=�/�)v���CaI�46��*� p��7�#�'�,*:�s[��>Z@�֦�l6��8�ɖ�8�b��/#<��W���ɨ�FN3L�4
H�	���Դ��Í&����'���6_��9jƱp�w��;��:z�9��/ d����卧�z2[���hF�D1Fy����8�s~��5-��(�ͷI�*X?T��q=���aɫ,QV_��g3R�=NQ���Q��;��мX7�r\еL�Q��7xҁ����Ck[���$�Qb�Fw$�Bb.?ͮ�bntje���:��>�'�[[���¤�� �`[�&#�.7���|����3����S�!1O����+���;�j���C���d(�����;�c�\��:�bh8l0��?މ	_5�����n�O`���O��fH���.vE:e7���<�����|�p|�`�����A[&��#|�w~sq�M^p(�r�d���b�&k��1���,��*67m��Ҙ�*���p�U�����������cs���� K�����OPB�:c����Cŕ��������r3?"l���5�,�֟L�a��h<��j<f��@Hd�s���,���9�¡@{��l���w���C,E�&�?}�HA��o}� h�t@x
l&B�����o�����������nt���a1=	k�d�5���inS�9��XT��Z]���@n7u��G��X����=s��5�*c�)�Y�5��O��NN��a�V#`�8��蔶H�1�x}̗p����%�ϧ�%9f�Sh6f1��#��)jh}��ፏ�ʖC�|9VS�f	}R�H���������Pi�>B��M�ޙ�7'���ux����2�	B�ڗ��OBڳ;ܺVP���!���Oq�mgts��dne�_�U5d0(��nU����EXFIIP
�A'�k�r�(?����ʋ�$������H����gٕ�����h���=����2�	�pȁ�4�
�e���t�^�V���orS-�\�16���N�PT1��B_l����K�1������uP9�`�.�{��u�ی;w�ume�I�����l�&P�!.k�x���~7���#��uC�c��>>E�u�ѻW�t�D�& �<_��ٌDs�m%��+v&�c��)�X� ���XS�Jp����0�	���v1�H��T%�����;��s����zb��ay�֨ ח��ت=�z	�C�)��~��єcU�D~;XF���넡���W	XW�jJ�0����!0K����k4}ْ%��J��ǽW�ߛe�d��������aQ�oe5��8`���)�%�Qa%.�L}��8��x�#��y��qZN�㛴`����ٟ;
c}�l=g�7O�^h�m�`Z�y��nP�v�I�\2��:��#=�	�Ԛf�G�6�y5�yL�Mr�*0�5���mŇ�?�An$5�|��t���O��[�g(5�=�,pV�:)�ia�h�'k�c��g;P�3����Ȇ6Ne�+���3�#rR�����yY�p�8�؛åi�O4��jV!~������M�)�Q{W鯂�渦�5j'�a������;ܭ��aHMD���e��]���S�Y�T���Q%���h2������HE��顴Y��U�s$��I' ���(��	V��w�*h��6A ����W�'ipDB����W����i{�8"]!M|���Q<�k���*B�丞��Mz^����I�13��������&}Ԙi>1�oڪZi#[S�N���3��e��C�T`#��h���
j�fH����~�1�1?��a�T5����1����{�"�Gv�Ϲ5�ş�s�W��S���c���퓛! �I��ķ�~��;���d-��Ál��RQ`5�	��|�E��YҴ2��&�2��M'��<�,���p�7�9��(���|*�R)q�q������&V5�h���q`ey�O�_�Q�?)�rw��l'��z��r�f�Π.�$3e���0b���m��r��HӾ�|��Q�q��r��_j��Ō!-���78y��l=\`�,JZB��q��"��Bez��˘Pֶ5*�}7�]�``��z�,����$�r��Q�Ng�4)=S����Ru����~�Fu��U��'W@u?pM�U���#�����b��$��>R�G��Չ�䉤��),�[��
AvSC��Ń��K�q0餝ZRz떖���Cq�"&����	E`�+x��'���tf�9�r���ΘC�-z���6��&�}W~����u*j�4=���Jt!��-��4M���'����Zy2���� ��Vn< ��x-@ҵ��ջ8���
���?�T_-(�ǋfN~����W���fB��<��|W�f�oCN���>�����͖I��4�y%�=�2�;�*en&>p>����Q��ڮ���l����jV���e��BZe�%p#���R\���a ��	b4'�Y}��;�wd�r�]Im�ǟ���=�Ɏj]��QX ��W��ʊ��w�l
�o5 Ɣ�-	�ӰЁhb�6
��皶 �T��>�"�H��O��3�~���P����h#��x8��ʉЪ�Hyᅮ��wU�X�y�h��Hɽ�1�h@'�;����a�΢|��[.�1C�<OV�}���KϽ�
�f]c�5���	�0k��(V���W��_N�Wy�>���A��6�v����|8�qqV�j�<�(R���M@��}B�����؆�9Šp�6ؾd ��^,��}`H��D= @���P��N���d���Jq(��:R#�O�ӄK;p�F=��O�婢Y!��m�p��z�e:�L�㪕z�YShwQ,���V�5�k�<��=������k��^C���F0����ҙ�2^~
	��h�U5�X3�<��q�ȋy��X�<5`�K�:aD闇@(H�|�(U(��M$����a.�8�%�|����>M���1l��Mۙ����_���Q�!A.�iMZ��U�mpg5�̙��Lm�1U)�X����x`p�^�r3���@����i7���H��}й�[Q����\�UA��Ң���&�+"
ҷ�8~췷���Y�AqxDT��xӿTF��L�ZK�j�MU��i�ˮ�����������#`UP���k�e�hV�%֡�HK)��]�ە#cvA?�O��i=J���,�y����S Z����H_����(Ƶ��a��?����Zfe��'��/bD����|���M�p Z�^6��KoP���~�݊/N�z ���	��+1
���>�W�#�9�ţj����;����]��$5�c��5N�+d�)���d�0)�L{�9�Jbl��<�t�M`�|���c�K��cĽ�s��JR]��vӗ]�dZQ8�ϱ�nd�rQW�'�q��GU`[����^�[jH7�I&m�0e�.���Og��9��ßpX���g~?���5;��z�o���ѿ?��iH�Z���غ��c���Y�����ڠ��y��0?|>c��o�k]�q�E;��{ʔ�Wl��y�*�dh�\�.潚x��_��>�˥�%ƍ|dLs:(�b� K���o@��H
�3����F�������1RW��4��D�.Tz���Sc��L����
*�q�'g��."9��!�c��Q�Z8)ʿ�
�N#~��W-��?��L��q�g��A'�FA>�b&�ٴs�Y�Ja�S��yD�[���XR$�a���lE#�H�,�.sL�k�1%h8KF��,߯�B����^�HK�^S��pW=b]�Q��ً����,<PN�x����%�?G�����< �Fo�ゴYb�M��jޖ?wT���QE��T�ų�x9�پb����O�a{�����z5隢[���mI@ٸ4�̒FT�Qa����f�N��r?d���L������>�s������\"�)�'_);�և8�@��=-ė$�ָ�'���8��=�L �����]��m�'��f�v����u�鯺�X�������?s����{A���,�vl�̇������x��K&[��G�<���AA���Q~�e��|�8W�cK6h �o�:"Ui�4�<�t:��(�D������Z=��$4ib�w��$�O�~T�R9��nU~kf�å3��Q��������,�S�R�Đ���!�@�[�]k�z�:��]��ZtCoD�� ��9WnGW���������H���_gS?����-3�H�@���%7(0h&̔���<���H�87j�A�}�|9�����0����*N2�sEae��8���K�y\P#_o���v���T7dsx��^�(�]�B�8���ՏF�v�88[d NFz���YωD��k��+�P�#p�Ԇ�qȯu�8�M^`�_��bku�z�OU�5�2V@�qt
�{��T�޲�=�	���57���ဋC�P��,8�;@1��1���-���fYǶ��-�\7֌����0���T�>�}6��)�V0�Vȩ3�֯ ?��/|�U�#����d�]��!�ta����~֏M��dzﰭ·���ʩi��:K�)����9��'��&^M���h,��#�A"�� Rqe���reR�a�E
f��oEL�X�P)ή���d�K���S�_��IQ�w��d�̈� �5%��>�Im�w�{��&����} >غ��'��}���R���؃N�9�h��SD�M�%w��ē�2<ȣ���~^��ʮf�eV��mCr�5�o�߉���6S9�*�!��~'�O������(ȣd����n�&
�p��1���O�&� 	�0+Z. .^�����o	&%> 2���"�i�6�M�g��J��~���y�W�Q�L����_���\�]�R���s��r�`/BEQ��Fc�����f��4�I�!� L����\�\.���"��Xיd�X�(X?�Q��qc>���Y<�'-�QR��%�͜k(2�_c��+@�O/$��8y�?�uh���M��8>#x����N�����橚�ӥj�]�Q�>£P��*H7��Y=����)�s�H�A>aDF'�96�َ������3��H#����A����
�`.�<�/ MJ�8o������Ҥ�k���>JZ��|H��V�j��|��sl��������5� |�?
�,�]l`�5��7��Pƒ��n>�l��(�!K�B��W"Y���*�����q�5K�g���� �cK�nY�RN5�.A'\N~��U���
=崬���ۅeـQ��0��&ʕ�t��}��K;��/�~e@-b���t��/�ot��Va��	x�u`/��)O��!��NHs���Τ}�^cI|{e���`Ȏ2�nɠ��I_|�]��NCب�����;˃�i�|c�Ȏ'��]�/�l)�ic�8>Ń�[:�	[z%�����yaj:�n�S��1ǏUh��ͼ&�YC}5�\*�N��HL���TLs)����������Q��0���M���\�����b�΍��uM!��E6�a�b$�DT���-'%��6?�������Lh)?d�n��KO {�[%z���u@Lڢ�%]'og
���0�� -w
����ݺ���'8���w��y���V�J@�d!�3 zA�rEۘ����u�ө�F��Hzq��WZ�P� (�%2��n�Bt����H�o(ݿ�ƒ�o�޼��xQ��-�?KC�\4���8<M?XH��c)�O�t�U�ׂ�y�?x~�c�p5N����U��Į�	Ep"2x-a�h��� s���G S~�8��f��(���F�+��s�1D�v��/yr�r� X
K�Z�M.m5�N��W�>_X,�f��ސ8;4Օ����ݳ,EmN�N�e��)3#V�g�ƌ��AS�&uJ�ˍA����K�8)�O���J������b��=�Y�~n���i� 9-�B��#�h�<��~��xY�	8!~ή����G���*���b	s�$��+��k�4��_]d]�y)?����Ȟ����p?�M�z=5w���k�4�c���D+U�թ:5F/�5u�5?��s�!;��K���y����ֶ1͖�ÁĒJC{���
TPP-rݩ�g����m�c=7on�Û ���F�m'u*��J^���JG�I*�BɁ�֗`m�>��贍��s��6<��#ߪ���e�~/�^����&�����Jٰ�$P .�U�f�p���G�Hv
=kR������1}8s�(~���|dt����|��V�)th;�(P����T���E�	nЄ��$��Ϭ����_�$+���
�)���4���:CƁr����d�E�^v�!
��=����)M㪖�V���7����I"H}�x���a�k�YV��f��WB
E�L�qj;�C�:��߃}�?�Uo��TR�=OΛ�� .C�"����0��pUKX���0 (+��Oi��l��?��|y�T~8��&76mw�L�Xw�Iv|T��*�o�����w�]�H!�tҔ���Q���z&k3nT^h%;�O�9x- �:Vd�/L���j����EnD����d#d��i���!0'�e��{;�yat:�hLt�����"n�w���7$�&+���� �FX�J=F ���-o����b�K9A�|�*�%֘�Y_v��j��:s�z�Zj(ؖ��_}{�!�*��~E1v�N�,�9>⑖`�iy&&�����m(�_���+��2��?�e�uXU���:���]��ֹ�.��nR�,ʁ�v����3,�"�jڤD|���}�#��(RXfZ �����g8!�}g�6�<J,�8W#��E&aaj�� � �y����?���O�V���0h�l�
8Q�m��+u�>����&4V�\$R� n�H��v��W��2i#��^`c#G���}(���������Gdw��R�$�����U�`�k>�dV �[ �3ЖI�˚�C8���y�@O���8��CN�u�7XDsb"Xc,[_��f�/�,)�1ɷ©��AO�5҆�_� ]��mH��N��#m�Ə3ye�sn��e�إw!mY������u ˦A^�Ի*��G���@�;������`��i6�B�!px"�`Ŀ�w��p�<N�GJϻD�z6�K��F3�W���y�B�C��GԦ���/n;Fg�����z�� ��8-iP��֦æ��O�|i>$8�U@2*j��:�A�"���z�����C�QGnn�)�d��W�^��E�,|?��PpM���32I�geΊ�J���d�a�E`�Z~4K�,�����,c�Ƨ�:��"��Sl�8j=�e�ս��R����ONA������N�]���x�����G�[
$V�d��R4i����F١ N��!�\&{ή�� w%f7`^�u.I`Fm�s/� ��r�\�w쉑,�[�+ 
�,KR��Z������?�<�#Wof	�AYz�b�#k���i��"�iqZ�	�Ν��8f�<�ƚ�:$���XL7�0���	`�=�{������*�R����%q�I$�r.�bC>%L@fd�@�n�f�<g�&�󮈞�=��9��:�� ���;��+�e�w��N���dI�p<��i�����o�8o�&��FE�K�^8��,��P) d�������:KoΦ؛'�͹�J�A����)O�n�_?���$�6	<��ג��3C�Q�85x����ې�M[h4��4���#�O�$՞ؔ�"�F3x&�V�
cj�����|�o�s�
}� �q�R�C��`�F6�F����@`�k����w���!���Sަg�´|g4!e$��V}�@F���E���"z��>5�>�e�3Q�/�N�(�Ƙc���v�����j��EMTW����{��չ)[�%�^V��P��o�5hl�gڗ#M���N�=n�T��'jߊ��/��b�N��[��v[f6y�����H���A��
�*��3��� �������ha�LO� �f����J�)3��~o�+�];�Q�;m����d����1uy��ǋՔu�\`n��w��go���Z�2����h階�q�����p?�R�9��c8P�W5������m9��4X����=�gZ�E���a+��9uJgAuf���Z�MCZ�5�)��Q%��/�g��]�8�Ċ/"��d�! Fz����d�v��ߠ\��P�~)Pe�}G� ���,�̀�<<��qrӒŹ��|4�i6j���&�[R3}��zX�	=2��>��e�	x����t��sz��zTE���"����!�X�X�"��4q=����4ed�!�4Z��G��,_���]���ﳍ���3*�w0ؼ$��W{��Tm��6��Q�'���O�@�R�4�k�9�a�{[�[q)��?u�Z��)G�`.�3���1�{�3��VS@nԗ�k�{�11AnI{	,}w�� �ë����K����<D4�d����T��q������d�ֆ���gvCQ�R�/���*�s�g���p�4я�t����t>Q~n����Y������������G�"n��uUɫ��~߅�Pܚ,$F^�~�ژY�A?al�����	����3�I���鸱���h���sIf�\l�?U���w����J��8�#�z`p���TZ��y)µ��8ɓ��F�*�Z���{q�P�m�@�5�����]\�-x�RS�E�w2.j.��@y��x�������[ �<;N�h��[繖[+�eRB�9��:��_�7]͗�!�I��&q�i��>;���mxYod�s�>W���3���&�!�ˈa��H��Ͳ:��1��jW�	bꅤVg���k]q'zk!7-TL`Y(���_Tm���"ʱ�+���(�g����:SR��Z.W��X��k�rC��׀`l2�6'��+�5(�vO� �ɹ1�݆X��Sֈ����Ц�TM����=+(���L*�1J�ǷS�a�����&�CO÷S�R����Y-?��H��KW�Y�D��)��FT�{�f��*�(�ӛ�;"'�Εk�05rA�U��t�H���e��PK�t�{��+��}���V�E���|QR&�猱�w���u�2:��q#lt)���44�ꪏL���!�/n}]Xe�Q�e�s���h�K�sL�zVA�Ի纊:�H;�C�#�X�wr!/��	e׸�M��z)��9r�k.}�X#R�+�WpW\D]���M�����L��0"�������
=��XH�F�����g5�,�i��>�KKW�GR�SvR�i{3�9dA��w�+���5�w���9��U����P�[���ڲ���{������Hn��߇;�Wfʐ�9��X�Ɨ�:��mro
ˡ���X�\�ᅁT�AU+�T5�ӴD�/*�+/7��4�V��$�Q���ES�r����m��^����౸�-+������Q�C\)���̛�.��L��U��Ó�c3��V��B���/ �1��s�\?�����u����qꇈ�P�%q��������g���؂oE�#�g�dR�!'M, uxXrJ�/�1��8mی�T�U�TP����Ǎʢ��)��hk���lmd��ҋ�T����\���B�\����3�^��O<+>�Y8I�*v���e��X[�ќ��{n��Z3^&�J0a�{���Z��|�'ֹ�*���6�;/���زt\��9&f����9�=�m9��Ku��}.�"�Al��x��ñ}�<;�46챞O��ܵ4��+�k��6w�]���t��O���$�����q+����&G��5��h���� 8/�Ѳo9U@���@��@ԯ�f��\��0���`db����6��4�Td��	����*a^9�y�zϒ_�Zn�G�Xva��џJYߏ���PF#̇��F0�lT��f�o�y��0�q�-ɽC�?ۍ���H@�����~�ڿ.�=�Ī�_!�3�d"�7��y�[9�ȍ�4Or�ҝwrjMX��lUS�P��̸���:��q�d���.*>TO%8@��	ͷ^��R�7��8}Q����A�yO�p�}84vR9�0�U!�v������d��ٳ�1���U\,E�9�!�;�&'҂;��s 3��>�������<L?a���]C��E�>Xi��ը��w|�,�4�U"e_E_�AB����	8j�3�E6�A�k]̦�8�jV�5+C�n3����~L.��1k�/�o�H��9��n�8���>��C��>�~f�(���i�t�>%�R���U�ِq���'Z%"�Ҹ�:?��J>.�0 ��� ��tK�G|����p"+`�x��L��X��diUҋ+�ʜ~���X�z�lwQ�|9�l)�7��#��~��L�)�m��,���َ�"5���n4�0�F�,��!�5f�r���!ˬt1�w�Nl�th��q�U��K�"�����\0����X�'�)�d�#\b:H�d`4�f�_��IW�m�o�cM�g8�={��=a�w�K��G���]F��N��r�o��V�Q��o*!2ll��ۊt2�j\�����F3�B��D�������Z\�m��Ŝ�I�~�yaԸg�A]����jo���+7�����#G`�]`��G�y��J�jD^��V�+L�|�p�&oڍ(B������j
Jd\���<3�_ʄD� /�8�Ү��(�1�g�ٮ_� �p��mq쩅�8����=���Ֆ-G�����X9y S�~�*�CDV���#~��1�������~��'��l$a�v�K��g� �%w�Ɯ��������\�z�m��B\��=/
ˢM��JD�tw��e��5�j����3�{�T�O���|Pi
c]�9u�4v��xza�ʀ��y<Vc*]4^v���N��.�^��������֨u�m�⎸���.�c{6BJ�{Qc��^�l	u�Q<�~���� �N��!exY��?+�@���[�7ۥ��x�g����k�̟s S��zP3*z>�$�/ \���g|**K�`��M_GI�հ��K��ʪ��/��9�h� CI5�'g���-��G?�&3��V/4�̛����$2�FoR$��MͲkn����(ߊmᆀ��Z�����?��ә"�w��Q�S���Lg9Jqv(�Z��;]����̗ LV(�S i)=��_�\`
c������v*�q^�H�Esi��^��7��[H��^l o��.:�+/-Y 
�b�o]�$�g��ҡ��-�6-�d��uv�NfV)��r_�����Ѷ�S��o�3;��!,�
f����؉C�^��V=�/�B��!4�/B���0�6�%�+1���� w�Y�$�yX3���� wu�k穅_���b͋�Q�#�>�C��6��U���C�zHI>:�?ٵ茧�H��R�Ҽ��u��Ͳ7�v���	v�6$�b�����wo�<6�XGf7x��x/#L.CS��aD��"��5(۾�!�(�D{���`�)6�Dp�$�"lѶ�@hQ[O��v8#>�n^]��L��U�nu���Ik0;X��u���h1� e��t��e��v�L�r־�,[,�!˔�_ٽ������gq��
+`w�nrg%�Ҩm��5H�u3����P�f��-��ƎP��������aB6,��_��?˦�/L +����Ms[�Cw���*TOu�3�Q�Y���)�ľ`�g�	d�F�����s �/\5g�(��1����g���A�w� ������f=-�r?��fh�z;�Y�܃?`6��(��4��2�U�pP�Hu�
����,�-��`p��Ȩo�2��@5�tjPa3����oZ�u
p�䣨�b�v3(���V�d���C���k�g��$s���3�͉�w�P�����l��fd�}�I��{)�n[D`��x�<2�m�O��1G>���m<0�w~�L�_��db��GJY5W?���e=?R�e��	i"Tp���wjå�g�sV�<L�1���h̵�]�b���M�/�ݴ9���6M1epV�2�N�;{���x(���|0�J��3���ڞ�qaɢy�P�zM�.:��
��3	�����Ǖ�O�����ǐ���R���8�I��)j'�w����m��q�E����ֻ��b0-��b�M����4�C���_�-��0����0 �4`�;L4��g�~�g�zݙ�2�?=�������L�S��!}��޲��ǣ��.)�nPIj�j��3�炂���ӓ)�v�[�A��IE�F 0>i������oR�ȅL�����
��r�����D�|�L�zY&��Q�'`��ݔ�_w�B�-V����`��/?�%�݋��om�7�n�(�w~Z���� ���"�t�wڶ�]7߿T:�Kj�F���f���w�e��a.q��~,��f���x�U�m�X�ug�C���x��r�4IC�XV��_4D�� rp�3��������%]`�����
.\�2d��w�	[Ia�T|+�44�!"�ork[la���������C�Ao�P�dڊ���J��m?`b���R��+��*��ji��@=�E��WIw�64C@Y�k���g+3L�<�tC9F���2oB�X�����E���(���^e��b�{�"~D㌛e��N�7��
6�U�73np�¾L�������g�IN�m��'��n�x���n��2�5	��CG�&��,���?GD����\��WZ�0S6�t��m�[9~%@��5��s�E�2ľ�]�ǿߖ����>�����.^8CF��Ibq�B+Ρ�y�h��'<��O5�քh0��}z��q�?��ӑ�:���x{�� dµ{?�����ۚ�~A�t�U#@J�i�P΁PB5����������k�����9H�^��`Mt;S��x�%���I,�Y�RY����6K삃7�I����(��.h.b �<�]1r��*W>�D�:[a:'��۟�R� ��@�,�<]�)�����g�.m:��󳹽DEz.�1a-$��z��:^�W�B��X�8�^=9�c��-�rS�a��N!a�c�]	?��EU���&oz��  8�C���q����SĮTt3��}����q�R���5��B�c�܋gX}E���1�����Cخ$B���L�%�m�����-�{�M�5 v��R!��O]�h=��Y1{ wR�fLQDXo!R�� �=�7k�JP�V0p��,ս[T�|7_h�2'��W�;f6�ZO�m2iӏ��<��z��ǀ8���N��ex�+ˏ, H��.@U�J�����D�7���.i[���������M����j��O/g	<C�����ӔD���`^Jk� ?b�DĜ��{���sz�a�9v�hudb�9�� h�I�)iuVP�Ợ����j���������i�����h�obɡЇD�g;Y�����ր��l@>=G��V��ΟF��������J{�R{�?�2L,7Xղ�����1���SwE�N�o}MGq�)�#�#L'`'va��a	�B-�of�:Ψ����?Yk�!��l��G:����cX�E4}M����xX;F�(���%�R�K�;�6>���� �>aY�f�_��&nU5�R�vy^(�JUXWC�ݏ�=t<)X+��0i��K1�o����!"����w����n�x�\ۚ�+T�.c|�3�Ci�l;�{���\�?�Z:b�)�l��
&WgTљH��l��yp�{������)\���1�ly1�״52�׾���Zsq�����r�v��E��`�m�jm��<�l��z�'-��|���KI�@�È�jv����|�RFq� Wu�ϝ�҉���q��qo�4
���7���݆�ӥ��9C���@�]d�?�4ɐ˝k�֪����0�B؜o=K��3(޽�R����n"������=���������e��	eHWh����z�a������1ߵ*+�Z���X�U���aᏯ%(!6���{�7-~���V�4)� ��23�SR��Q%1�ٳ�8��R��FCJʖC���rۗ�"�>����̛�a<�����M�3�{zu�}o���)rB���'�+���2���qL� ��%T�`8��T��ϟna8��?��FN'�S*V1�fm9Q� N�i����Y��N�QV����.�£���G��R���։���	/�3x����g��;7��.�⥮Ǥ���7=I<-G�U��w�:�P�@�l���(t���ZO1��V�២i�ӳ�<�`\�/��W�R��N)���њ;��-��!�yM:����$�ڀJg�5�!�;6�K��A�0"��iP���N�Ȫ�����oe{�l� �����c3*ݪ&hխ�)�)XL}������p��VNDFơ�O�ͮ��
-x�uW,O5L6(��Z���e�t|��Ǳ���Z�����_p��g�FerJSVF�1_����)r7��pR���mJ�6ZӞFw@�n\������4F��g0nÞe'u��U�4"y�B�'�#N@��i�b�I��A7IsJ�ɋ�=��P���ϫ@�b�yј_Fv"E�����1�B>�2�%��).�n)���vd���恖 [/O����Z	����;,��ׅ˪��������VLУ�(�v݋���{��0����j�l���)m���O�z٦?�,,yXg������SN���DD�j���(Z����p���9r��{G:�V��f3/�]1��m�z�l�{�ѻ�F��RӼ[]��haST�b��t�`�����h�<eɣ��]���'V50�a�{��&�ޟ*m�T��^����@zb�����Ԧ݇m��;�lP�'�r?�LC��1�x�wK�P]^�d��E����O�B6P����.~��A���?/�͒�?�I�)���!-�2a�Ed?�;к|F:�Mn�\�����%x~i)1k��AA�L�\*��c���e��vW���m!���u� e�o��6��;f��Z�
�K�Q��D�U1�a�{��=�^��TJ�oOn
��|�4��� �����Z+$¢�njI�U�#ߔ�\45���2�oCV��7u	��4w@6�[�:1��ޏb�B�S�!���='쀮WD�Ny���?��gd�W���/���������@"`����#y��q^%V����^F�G�#Z}��p;`B#�
_z�S��`���R�����%!m��s�Ug��o ����6
������a|t��O��C�A�a��_Ew�V�<���pcP��J�$��
W����b��\�4���Rb�$ߍ�R�p��Բ�n^�_�V=}���CQ�U��V����{��ҧ;cG7��>e�~�׼�+�*+�y�b{�%;KE;�����9��V�m�Ry�)�l��R���颻`��C��2t��~]5��O<��2�z�%�m�,H���h`��_8��>~��	�[���C�˷DΎ�թK�ɿs~����1�Me����]	8�E�2B��Yxl�&�v�Zc�pexN7��ȋ��o�Q�+�&a.Ex�Vr܈r��a�Pu�L��S4��0�z�c2Ì��3W};²@ϧa4I���e�������L����f)���2�CB{��(�9�m̥�ɼ0� �\s�G��wʋR(�>��*_1�H��X�*�+�/-�.V/o�:U�gz���	�a�m"�%g�2~f��C������OT�cFV&8Dd:T��r�����S������J�*גY���KIJq���$��9tY=`���7�Q^��<��C����_��������P�?|���� Z8�8K��3�d�s"9 ѫ�q?Q~���Z���+y�����/o<� ����&fh?��K�"����
8]�������zC%���9�
�s�I���/ <s����q |]�T�Ҡ��:����^{Jcٵw,�kZ�L�φX��ӽ-���++˯�h��U��D��?<c	��q"~`�c~%ׅ�"�Q������ro�I�_�z�&J�����%��'O1t��~���;}7��V/��3(\�a�)�\8o�qO�v���d����E��e!+�:q0yQ|�\:O^�����K��`�5���=8���� nh���lƏ��b좄�Mx��c<q>�W�9�wѢ1�3�L���X�1g[�MJe���(���V�TWd��*�U��F[��7Co�YV��~���Ô��=�8&���A]_����B�Ͷc��H�9���.�j�\�83�M|x�Gѭ���������ȵ�u�(s)8H�|:�j`�<4�<h;����*��L��Qˍ��Xn�ه�՜��S���G߇OАߌˉ��΁ג���ڵ8<��oU�˽��;�n�T/��9H���B�ޯ���gW�������"��+�!�5��v����&�[�d6�fz=��3;��/�G�)�sD���Qop�	�6�U��^�l2���%bR�/X�:f��Y_EY��@W���Ű�!x)�)��77J"��4���ȇu
~�R�φP�3����$�����U��gn'���S�u9�m�VL����2�]f�����K6���
u�{��"�y$O��~Z�C#ߩX|o�����_�aOl�u_<���`��vLܛ�~��w:����#���Z2vu��q��\��k]��l|e����2Wr��/,�"1 ?n\��^�a���Yhjg_ϳ���+.��j'�ZD$>�Ґ^x�C�d����%f��� ���| �<���3v��!Ţ��kb�bXr�Nr�:"�,B�t=�
@��+{�_�*�=M�Y�{<�A�3'�`������0���!xZ��s�02��>��%A.s������
50_{\�����MN�,�9����|�u���y'���70mT��R_�5a�2�w�1ʂ\^`Y��=H�9�f�����o�F��n�j��\�(`��0�bEʼ�+�²Z�R�呓@�Do���*p��T
����B�\h-z����+I0%B��U�0fM!�uŸʀ�U3)d�֪��AaO�#W9�-T<��;�^߽�A$HxE�btk��������~7��x X9��+�M�G�_fx��m�L��.|�ea>���i]�R�o�k(�$Az�l���n0�~�݆jt��Ke5wZ ���T�M�0��j�9vD���2���r��lmf�܁9 �B��PT̉����7T�����d�$ ��ו�7��5�������h_�И�mج�� I�B�D���}���ך���a$�
zMzY�ejXJ��=U�,���� I?��(�_o��]|T��Ey~q84G��F^�p�r�a���"��.F���E ���oSͻ���L��h���6�x�Ԫ����m��P,)�\1mی��jr��a#��g p�<�1��F��m��2�G5�q	�@
eĈ�	��~K���7m���x�6�Ë��{R7��Q�	 W����[�M��,[!��Re	gXd1Bif}m8|ַe��\�w[��!�΄
��9S@+5�Zd���G'НY��̹0۠m�J�8��@́a���r��i��֣#�rh���K��o#m���RS�r�eXO�Om�(�w�r�ik��q�b�G�Dm�	����gZ��|;m�~C
`�ML/�6΀s��4$��E�������^�0��ـ�Z��λ�k� b{��繓�;�UlRÞ��� �ԑ�L� �B�1Ä�q,֮l�����������-<�)��4�kt��P�n#	n�����+���A�ި.K�%�6p$a�8��wAe�x4$��a�Z^F˒ݒx6�Y0@|�٧U-7-��ֈKb���`G��Tԯ�F@N�nt[�"d�_]D�6��x��
B<*�Aa��߮�����;����)�\rd$d�H�t[wPJ�������9�VTş.VC��91Ń�WED���d�C��e������ۘ��?`[^�p����ф+b�AY�$��6xp���@?zK��Q�|x����Y�I��%'X�ˊBԿӔ�{u"r���W=y��Z��{>�z9�$>֮)� ��'x:
�|/IK�T��*M������D�����}�݆���Ӗ�c+b�d�Z]QUA�)X(�Wi���k3��87En�?�+{�H�<� �V�g�ۑƖ^B�B($�䑻R���KS�e;!`ps�e��t$�٥b*)'N��B�%u.XYi��✴0�Eʌ��<��O^��7�Ԗ�6ٱr���>T��m����3��(k�4�/����F�%;��%Y�:�����Z���Pf�l�V=�īiV���Z��af�,�����4TdwD�%W�<�s�蟎�뀪D�
M�����6,/2��h.�����<h'#�,`�����C��AU0@g�Y��nEZ$c!��'|锣3�dDv<��Wq�������u?'����J��X�u��vC{�oL���D��ٙ'�������BZ�T�[�dC�j��jb��]>N�9�T\ԓ�)NV�r��x|�Bj�%8?<���	��U�,�ّ$��Ƙb�hu��)��d��t>,���mś�܉eCH�l'�ǻZrܞ�9���~W�Ǐ(��{���v>�9������l!�����Q;�ˊQ�*�����6�K��K���<0qs�����&dM!Q����~\��t�VN���f�H?�5�2��p���l�_9�JW�}��'����N���:�[�܃MLDx�Vh��G8�~�����w�;������U
Z4V��ʵ�����n��9b� ��),U����C��E�f���&�h�:��#Xc���mC���~!�g6Ӡ�z��O��ˣ^��'��\ʸ�1��q���q�,r:�5]�W,В���I��?�=��L�_tf����2��*Q�����F�'�{*]W>N/Ͽ�)����2��Z}� W|lA�\n�Y���'2'��F��6�~=���wb���>�M�Y�\<Б2Nȗ3I]�Cݥ�2�Ѽ�I���W�® ;��َv�f3��"|Kx]�T�ܼǜ֗`WC'+�i�d�Pb=�����D���X�����E��g�J4,�H; �����8+̐�q��h���W�hI�����b���g�2�8�T��_�p�]`�F�`��z���$�c.(�zUA�n6�	�0#z���1����p�X��G�Ec˅�R�҇<�T<��C<�+������y5o��d�v���S���Y��v䳆�U��R��~�gQv�γ<͑�"Y��CEN�V6�0՜�nT8ȜS�
�J��|�iS�ctaA��@�c<��!k��?�o7.h8p��RE�Q�BLj��{|����\G�9Y��X}XJ�d&�~�6�q���	��Ԫ'��чk�Q�=�Q[�D;�"G&�+���^�˼��?��ed>�o̫֝
|0 $M"��I��P���B��	�qH	��fy{s��nu�?$���� ��U����}m��3w�ĭ]�|O;@�����ݷ=�dI��	و�t��4��\9_��	<��d��kA,s�?n�Z�
��w�۵��L��Kt��|�h�5_R���"6��R��0�!���|�k�ㅚ�YQ�����h��.y(B�8ä-��i�1r��X������	�j���:k��>ɛ�pJ�R���n�J�$1~�[�v	.�G@r��~ir]����%��3����B7��lɆ���0� �]�$���rE[��]��e�ˤ�N�b���<��f����m���o�rDN/#��3߀��䙏
J�߱���Q#��w�.���H�n E������4��d�o�Na�[�yw�:P]���P�P-p*�>�W$�%`��<	e~�aE�k�=�:FBO#i��V$ÿ>I�[�1�"�g1������g���f����Å�dp�7�]x̭��G'$�ώ��pnw���){H=v���`���+������9�F�1�K�D$�����M�pn���$[sV�ȿ^�����@��\N|���|�R�91M�v'j���Pg�.PC�`�!�.�_�@s|ٔ�7=���s������y��p�D�/Ig�������/�0�apK�e�.��{%Ε*Ҩ�&-��K(����.�eY���'�d���	��.�M3h]����&�NW�&�c��|"&�4Xl�W)Mp, ��uk��|���N�E�B�[,Ұ����#�Z���\�������뇊;�~�]Wv���� 9�L�$+����h�薻�>ys��7iӶ����=6�'����z��s@?�EQ�>��o�c�
Y��"*�/�aJ;u[��mBT.�u�W6�;��K�ݿ++٫:��v�|LW�D�� �Q���0:?cG������f ��?&���5`��c�ɓ`|Z��j��4KxSَq�zf���.�;�o��j�]2�$V��aX��W����Nu8��4P�!�E�^�s��0q�^)�;�%
Ae�+?3���H�[eG�����2o@`f�nH�&�j4�$,8��Wdzf�����"x�6X������H��5o8q\�IY8(
u��/�S��Ũ��k����я���f������~�g���%��`�Pҷ���,0�~1oY��c�y���{
$m)��/z�y���2���+1x5K�����F��!�}r�Y��>�B���f����_ʿ��d՘C$dޮ@�L�Q��NctZ�u��~�i��5Z�R����]!.W�!��Wh��Ǜ�6wO�f���������1mu�x��*��hY���J�M�����c�7(ْ	#s����R�+���^	��`�_�O��+QWM�j��V��7���^w����q�F����a����T�m+�������kU.{���_�L�Sܩ��T�v�`�+�ڍ��u�ϸ(c1�=%y��f�${�U�)T/y�І�6r[54`���?q/�m_<Ac��:��[
��u'�eg?�:Z,��&� �N�2��W�5j\^cb�������m@�� @�=.b�\�=�=mTÜ�I^�EA��{�z�_�A��ŶM��9�|�?�:T��_�<|x�� >J9�d~�j8��p�(ǟ���^�n�{a!	ȧ����)g�{O%�%X�)u��iu�z���\���b&y=��j.�q�R���k����Y}���x���c����V�f�D�9`V$��6�2S �N��3�/h��4�����E~.��~o�$��A4���32�Z0Z���[{1�?��:��)���w��3�w�	�y�-E�8�|Ns<vg=\b�4�2�쏯j�i����� ����v���ʎLy�HEl?l����l/L�~G��U#���ɯ;2o�U&m�%��=���twak�_��� �c;$Nw-��:XUƮ�s�DY�/����*3qB��6Y�M��[�y��I5U03-$�\��æ��38=J����|	W�t�T�D�`C�\B�)d�6^7��v�h^�N_	���m[I��X�O�o�v �9��k�����L�o��z���¼rӖ�!�w�� A��R�RN�
�sx�ܵ�E����ْm��o�'x�k@����p����.2��㸦�~]���XY�A����K��Dx�7������v�xi	K�j}?������mT����>�����G,<	�(d\��]Uk���&�CQ�ED1f�cK7O'�P�)q����	+���s_���?X��DʞT�v���W���Z�:A=���F�M�K�)i ���M��,�|%@�Sv����dJ����i^���jC/j@���b�ݙ�J�p�g7u碙�#@w��(挂��ҝ7���%�8$��o�:�bg���sL6�� =g��&�72����������n�D��-+��"Aw7r�`i�g��f�:ù�o�Z|�a�=1zG�p��䯾!�:��e�\���A�q��!�3�QO�-����M�!��>$�G�6�{��x�WUH��O�S��_Q�"����^ؗ�1,y�O���h��!NG�s"� Hf��b�)�#�����˦���dX����_xf��w�̺����l�P��i�'�\r�VYz����5>�5Y�k�lp<U�#EA���L�s��l�]���@l�>�.q>i����NH��e=��U�o�M&u#�8?;Cba��<!2�7+�ehb6.f�aB9�4�r�+ĕ��*C���z
��ۂ��������Ϭ�<�ک,�n�����e�z�����CJ��-���2��;��C�.�<�N=�~���W�����S�5yIO��Kގ�2`�����|��#���E�TC�M�t�o�U�f�<uV��	�����(��=��4Ղ�lE�ze����a6b/�O��O.����[R�T�z�U�3|O.������d���%�=ֳ�U�M��:4�V݁`�_�&
3�?A�����@
�����暈qt�F���Q��u7y	�28T7�#CD<�T��wJ>�o���ge��<��~���7��|��C�#/����E������W�&��{0 a��K*]l­�#?���;@��"3��(�~�1z*&��7�����������Iẋ	��&�Z������D�"K?�=�׾�Z��3�#����Y�ʁE�Q|<�X���%�|e��I�
 �Hq]�^-�'ӵY��M+ ���w��Q���P�i��(*�(z�h�_{[�����0��ޓKid�egN�}����n}�A�q��$I[G�V׀9��W�L|$��E�앱P_s��za��%˸�KO�B����߄� �<���[]0GT�umm4Ԕ�j`�@�R��Ln�{$����0a��	1����H��N��$������ԍ^� M�ÒLP*�<?����x!3�u�E�O~93��bYۂ���(k�55��dQ��X���ϫ�Pf�<�N���B�,AB��
%G�^!a�a;-);1��@7~�)6��-������z䓺c|,��B�q�t�I5��̍���p�[�����w�\b�^��k�J/��)t�q��^-���"������KS\��^O�Ä?�l�c/c�=Ou�e�M�=��d����׆��!ͿYk�##�=�To�e�#" #l�AY�����W~�ۍ;y���ZI������<����iˏ���͉��dN8�VFl�����l��J��5(x"��9J���p��f��f�a9�Ja��we�����*�����jM�ȱ��?O:��\�idWdn�I|Ѡ�O���W���VC&�m���	oZ_s��4�h}f@j�u�R���Dai�M��0L�"��#$k�����F�%,���`lf����pZz}2�=���i�ƙ�l�VS�ki�a*���{���Ǽu
Q�:ɟ���5t3�F����$�[r �X�|d_y�S�iu����:s�o��+��G�2��}&�i����I��}���pRs�#V�%�`/�(���y��m�U�+4��2tɯ]v�Q�O)g�a�_�m.;����w���^�6�Ʉ����>�c�Ov�1y���Y	�ݧ�j��ݮ��mX���Zh�[�V�_͑t�S\1�{)wv�2Y-3�F	� F-zc�6B3aΝ\8|��ݯ8�!�YN��M&f�.�?���k9��@��(J�|���-�֜��f�]l���R��)���d��Z��c�k��󭒏k��sQ{w�Ǐ[ۻ.%V�ӕXaF)����-�6�q���y����a�1�� _�U�L]���S�
#���q�q~Z�D{��]	D���k�QK�8�q�\�4�����}IP����X���^��R_� ��b�}5y���nr�ee�,�u��}Θ�9ę ]�����ȭ�4Rt����oD�Y9.��}��.9�%~ד�z$�{�n��͹x�|�D�����=®n�-~��B���Q��\Y�:�ݐ@�vb����r�%�<vs��;?�ۍ����@ˊ�`t7{���A�7�+�f�,��
����3��P��[��ep
7܆Umq�4nBr�,5���l[��QR7
�����>xy���ɋ�K�FE�jac{���C�w1^��s��M BG�EJA�2��`sQX��j͏�cJ�������"e�]��r1��$�z�ꤡ*2K��n�E$b)�3�/.P{%�|�FCFG��k��]���#ɇ�;7^W��?)�~:�L�/*{���^�?6�敺���+p�Q��f8���Vha����g\�	пc���U����)[��Q�;邚��)ň���� ���� b�	���V%�����Z7�� �,q�B�3����IЙ�S��=�d/6�O��`7��H|k>�7vA��(7����z��`��!9rH�D3�]���$��g�^͋����-s9)K.�[E5XV�4$�b��v֥_���c%PU��6��sYџ5���ŧc	�2߭d6�z�}ilL�`m���1vrq��!�5���~s\�?qU��[bn�Q[j)�=���P"ӊ���]db:{��S��L��f��@
�<���a��Rj�P��[��3���W)��|O+j�:+%���'�gŤ&�������|�v����B˼J�N��-E�;$�`A��q�ŧ�#}�T�-6�*�C��7��e�%�ۯc|�"�
O)W�����nn�Yv����Mk+NX�>_y�i/�Ɯs�3;���,��):��!���FjԤ��kvy��0�(����(�.��K������,C��4��i�1u�#+�$�J"!�M��x�dӽ���u�m:�n��tc��ߑ6oT��""��$ֱ��Zj�MAA�˻��\�G��0�r��o+ �(�Sz+Y�e'��C�,�[C���9�S�Z�
�J^.b����:�1dw���������2nE�.+S։��!/;�$%�?ƭt��[��psR�R�TH�V1KDj-tZB����u�#Nv���6�A2|��r������V��i��(�+E��Pѧ2�)��!]Va�lMP��|v��0]y���h�����&�ȋL`"�&�@���r������u�h��q�0Ni!m���{�̂9ED\�O�6AZ^�sƊH��+��q�dN�O�����};7�AsI���]�-�h���BR
i�[�Z8��:)���`@A������Bg4�\�ʗr���jOz�}��6P��g�jB�r��c�#sd��B#fҥ['�H�P�,$�����!c�AwcN�H� E�(�o���F[��ռ�84�oݩ��jQ����|mS�]:���!�x�p�_��E���4dN�8�@v6�ʶ[��e�R1�K&�C$����#�A:����H�h�ѻRn����r�	v��P7��$U#	�<z�z�b& �3�--zG�W8 �kk�8�ŉl�񅵞��m.����Y'Ŭ�f� (d��1���
�eLP��
�|j�u�ܱ��Y�IB�����$�u�2�+�}^~]d@;��� <w Um�k}J�Y�b��A,n���G�ŷy%{�e_ y��p�;r	�)���^��ZvDB��h������gM%Z�U�1�J�1J{Gsv�;�!�	w�U�N���m��4���U��3�Z�VI�U�wO,_�=!�g |��âDr b�,&�2HN.�� _��+s~;e��K��3ϰ�8�9��������,&>�Pﻦ5�[�&$1{����>��A�	w���n��%V��D�e��~M#]�n�w@=�㖘�6TN���쬽_@�8=�7.k.ae�xI���ca��`� "F��:V[1.�a���A������c�>h6q--���7���pɀ.�^���6"n\�U��
h�+z��ꇚ��Wl[�.H��( ڰ�S�ء�fV�,���0�+Ի��`܃�(�E��*l�Vd�7�c��Ԁ�VCǞ�$�;R�2�W{����Mt����ލ��u�����H�A�A��G\$��~���aV����鸎b�>�z�Ge���u!����,�[7I(lq1�;Q"-�$�������<��R;G:O6��F��H]r�;-�1����� 3��C�>�.�hF�Ks�^���\��H0a�Hሃӓ�J�>����2�+EV�C0B�g�P��R8��!,b�I�"OZ�ˉ���ؗ�e7^��Ӕ��C�`  �5c"�f�[{��V:@�$�0��f��⯡�zՈ� }�,�.��x.x�\��o��TY�Ykf�|% k�p%S�l���a��������KAN�0;;jj9T�f͟��w���V��B���|/t# ��Mk�(�E�<�*�����j�2�/��7~I��Q0��1׮'L;gT�g�F�=�ܐ5(��x�-�!���#&�i���R��0P����� ���l���6�[ �E��}��ފ-䲵V:����+>���yG\��u��b�;��֨[5�O@�E��f!|�
FL����m�a���z1Zm�NUZw^��<#:p�Exdt� J�I�yŔ��n�&�99�.�[�w�����ݞ��J,��z̚�Y���/?��B�A�=߂gs��q��`o�;Qh�9rǀ2������7��o���0�����s���<Ɇ�&og�Cw_5U�uQ��h���1�蘒nޣ!`�I���YJ��OD D�!�Q���0���t��;����w���81��5�Ҧ�R���v����)T;�6��^.�iջ��9��+���2�<�8Q*�K�CF�2~m�~��P�Ft]f[^��|`>�/�<��N����������u�*�F�#IsE��1��,��%\�-tt%g�I���3?�n>�F]����Y����n̛��0K8�]_E�V��F������u�N����=��&9�w}����q�m��X�0�)f͐��Q����A�h���_X���%?3W��y����O��o�VU��ɠb4>?�ug����}0Z�3U��e<W!�##�:~�)&�����j������|¸
���a�'8T�s��Q����ȏ���F���̯{u3-Q�`C_9�V�K� 9�M' �ϳ9w%�$������2�}j��Rk��Z�Q\$*u5�ǲ�sm)�j6W�7ϫ��T!��,$2�����ڞ��P�})�]�t�i��|w����}�$$Kcpo� �������6hSs�S]�թ��HVE��}\N�lS%c�p��~�w���Ȯ��$F�!߀�f�:툉qB��
ȅ_��g���T7u7���'b���K����A]���Հ7������H��?��|`{J�/ЋT �Vӣ��������u��(�
�S����aw�y�+x8@{+;����0x,�R<��/8� �J�w�����[K��YQ�q"�u����u"$��w���Iv��I�7Gj�b�<�w����'�G}D�U�+o�ZN���u䡤)�����H(u<Qm^��4E�'���5�9z�����h_7�nA�C�y��Q=�����`w_�O�l%s�������^�� 1�w|wm`�w�j�I�z��TԮ鹽ǽ&�h�^�Z`�H���#,�ت(=(Y[rvZ��Q�}��x@=�?���M{���$��m�~'��R-x�l��0���W|����״pK6m�}Q�Fϻ��I0w�|����>Y�P��Z%���$L�'���q�P�`,)IC/*��b�JE��*�ɡ��힓J+�����F��#�$esX��t��n>\J�
���|o�9B��҉�@�����L��r�y���8/%���kiW?��(vX���M�BZ���HI�N>�m6�>����fͼ�ѿ*E���'�]m�y;�A�ּ������m�?7!�ȡ�B����$�T�z	�W���(�6��o��t�6�Ƒɡm�*�D2�^��Y�v���:غA�<�����w#M����2J:(TfP���r��%2�%i��2c��R��|蹾-yC1�20i��_4����!�+c�T����ۛ�W�!8�)?_vȕZM�P�ӔKKR?����n��?N&�9/hu%�XjB���'Ñ����93(+���c��_#���_�nH��¶^Zhb�i��6�7m�\3�|����T�J��n��'�����.)T�O��V9�WX�\���`���'x�^".4}h�Y��oz7-���v�ɀa$��kqĆa�k������у۴Nְg�TZ)p�; %`� !:�g]4��;��ηk�&p�xZ��̀	���8�s����WFd����q�_ �F%��KY �Q�H��N�������m����y�����	pN�h��<�m���Ÿ��	��F�d�D6c�����c����Q&X�Fo>`��={��7����A�b,ه�~Fh�k����vv}|9�9ܝ�rE�|G�Ԏx`��W�ݰ;ci���p��~|PI����h���X�i)�����K7 	���u����6*3�a+|*��J^te��z"	�>�?��2ǃF>���f�F;ҹ�(�u�[����^5����m��������a�-X�I,�CBO*�d��gk��Z_��l��f�4�8�G�|��݉%Ѯ/�?����IӃ�s�����vX��{`t>�z�b��A6m���}Z�䈮%r�7ۓa �%��~�(W����� �Tfvۏn�NI���՝Y�8׳��h�9���5��C�K������<S�ϋ��ТE"�c_-�n�U�`���2YB�s\��Ɓ���a���^�FJ���Uk���g�V@�y[�^^-Ŝz�x��Q�a��#?�;]�%��xf���N�<H�U
�6!����D��k6-���]����vѕ��t2�O
pi��{��Nc��^lBϹY��p�U:��V ��
AC���<�[�u #�6%�j�<�wN�]@d�Q�"Lzs�j�!>@�������t?��9@5��&#6)"�pS����Hʭ����R"F����3u��Ĭv˞%��gj��ōƮ ;�;f�㏙���=ul�����`��.=H���=�e5�z�(9��{g<s?�eئ�s)��6��~��w;^"ʻ��"&aQ�S��.N�J����9K�����-�����L����/E��V�q�@/�l�W��Qd���llKM�deov6}�"x%���ʥ�7�E)Y<�I���ښ?Fv桧���°P�ze�5>�ٴV�>�Z4NEn~���pa%X�l  '�����)}� �!Fry�!RT��
�Z�����,�*xа�n�|����`������&���Dˎ���o�h�\y6)�Qp$-�ؔb�ѯzz��,h_+�q�����?����u@�A�r����N̜����D�:\oΌom�|4����X��`fM}��-�YY|�3-�5� 4���G�2(�lh}W��I�ȷW�_��2�SR� ����VQ]Q�dAޘv�i�z�j�1k�u%�����S'b�ysB�1d3�B�X���Y��đI�~��!���▙@���.L�Ry��'�A���p�F��wǦ�F��LbBa��ʷ4��Fv2�Μe\W����-U�Eo�:�S�ᎎ��U�:���u8��<w��|-�g�݇�떕L)c(d���hR����ʅr?�����P�n��"�ا�%G��u����D��%S��*T���f)	A��:�I�C8R`�2f�u��8��Z���[~d��eIUiıp�<[�K�ŷ���zsg���AV>L�Q����N�R��߈A(��	����BDP+%#^��F۵{Ӵ��I��0ґ0?��&��r�P�����o�(���^H���#���oη����/g�}_�W��
�ua ���h��(�oQ1��JL������&�Q�����""�5L���~��C�d���M� A*�?p�h���w�̿},�m�V�=*�(Y��,����p����].�B��g���νy��	��F��nV�1��ZѸ�c<G�D"NX4[ޠ�b:�<z��Y�Ӑ<�����5�	8�Hz���]�0��f}�x��K�?��q=ԓ��5?_�O�W	�u�CM	�A�������Z>��@v����7G��!6EBM�}�N��npi��n��G˅����VҦi>_l�^��.s �"�\x8@n��<S��屟&�_i�r��n"���g��Q|���0j�`i�<,���
��s��\�b��$���-r%1$��]~� �Ow��Y`�{h1)-f�.�̽�����?R��o,�x�3+�������П���W-�2�kW�T2��4չ)0�<!L8����i4w?���C�L?�7����zU�d���53�la�lxa)�	H?|�4��=���\�����Z�U�3b\9l��#4$
��Z8�H⺞�q���5���s�q�����== v��+��RS��3�Vm���!w"�����猾:(��"8�v#�ҜaI8�j�U/�Y.sk��� ���o-�O���7s��z
���g���]��D������⓺���҃�y��Zꁼ�W�>]����Qy��`�Gl� '�-m)XXeBx�'p%*�|�{�D�p�RyJ���f���������)���{��}u��g;b�_,��kX�	����h�W���xb��?��-Oa�6CNkJ0�	bjش�V��C�9�p�I쩠�,��W�EMC�<���GO	�S����o���5/���ļ�p!��wU�^Ry���<���u��&19�j�l����n�^qH�zoi0G�>4C��"]6�KvG�����v�*�����	Un�
�$�A�$'T;sF�Eϒ?li���V?/���*I�Q~_����2��ږ�uC��r��t@���SM����(����:3@�߶�{�y&-�o����3fS]'�/cXղdc�*��O���?Y�#�<K�Q��H�����^�'����d@ ��!����b%mt���W��c�U�Nh���g+g3A�g���UXg�����]�����n��}a�<�X��o[��� o�0K~��$�s���=|FOV/��6|]wD��X Ӑ)p�jO���jau�+��>�w��%1e���$�p��G�!��YW�f��j���McH�$Z{vۄ�W]چ�I���I��������~�C���WSU�b��,��	�|�ߡ(:&m�s˅��r���pt��
�6v{_x+�6�4��|y3�?���C>��-h�-�NSNb��'�ԥV<��x"��3׮Ɍ�@A[��+7G�J�Yʇ���+����Wk��S�X���4�d-��w��* p�)p���|�+��i�y�8I�0r�yTֲ�2���i7����9���d��c��ɒH-�/l&�3*�.f8G�f
�<���;%�A�Tm�,Co�K	Mן�s�D���5�#Y�dP��:R���y�T�d.��Zցea�;á���-0Q=�z�|$F =Efw�lV��I��b�c�ǥiT2b�S!�4��+9��\���� E0��n]���/Q���"�^fy�n�@JuǃI��!�Q`�~ h|�e|<2��������E[�E�_���@�N�]c}c����]M�O��<_5�ځ���y���W�]�Yl����;��_���S5�e�w����9t�#9��w���f��V��ES��._��|cpڃ�f&�s ���W��:�ԈМ�		�iX2oOW?#��q������~E2�b%P�ʹ�b�Nj���
?���t5�h!X"3�Ӿ9Px� ]���Z��g��ـ������݈bl�^]޸� g�k5c��X#U�B��������h��W�)�͋o��o{c��~Kh"O�y�Hc�I����8+��i�=���k7hDr
��Tz�Ma�K��b��� t��}s1����$���EU	M���Ou ���M�K|��G�(��v:�+������O�c�v���
�G�q����(ԂM�9��y8Ts2+ 3���g� ij��N�I��� "�S���ian�%yO@��*�m�G�(��u޼��H�1S�0�fƳ�{s�&� �|�]}�O!SNC��.��WÛN��B-`���Ǩ��G��[�TOq�\��`�����?��z��A���rf��Ybe�����?�PC�=P;�Ü�3@��yƆfz�2W�(��9if�p���y��[��T�n�R_I,��N�>)�?�~Nۋ$"QP�Ճa�G�)ДN��(����C��,�ИA��+(;��EL�����X�s�}�8H9C�.M�uN��1y?"sz�tM�N�¸IN��HA����L�n�3k�Ua���5����4�)���
�z���_��dM����0�A�o��6s@��<ϰyx�b����_�F��>�'�~�����"z׻Xqi��?B^E��<"��u���V�E�J�=��<���W�EK;�M(�$bI�(舎I!�XF���-�U�s�3w
�M�Ny&D�k+Z�59;���x�/�"Fe�D��� �.��`Ƙ������8r�j�oߋ�١��t��)B��Sy;n�?�2�#I� ��7	}���y[��*－ϭfK;����^"���{S��V��4u2�!ug�7��H�J���6����P2��l����t����a�{֋4��������cOD]�(B��(�!���#e
�6J������I�����@�X:Y�����O� ��O6�qų5]Ԃyj֬ˀ�[��tY�+*�/�U�X�c�-f�\� M���l�`������?>��On
@A�M�Dx�V}XB�cOGL�{w��v�z)4i�6�!�Gmh��$�N$թV���1�w&�++�({S]��=�����G�JA���:��):&A�����$�&���fm%�r�����&���\��]�����L	o�TO@t��i��d�g$B۟�}8m�B�_��{%��-���53������v��^y~;^�A<{��xl$M�ʐ�#�Y���(zUY�y�E/%�H�ʢ�����!\�xB�VLʼ�wy� =�0T{?k�8��Tq��b*Wl�Sa�#<Ŋ0BV<Ǵ��C6q{ ���P��n�6���9�"�s�3�����)�N��4bV��_ڥ��C2�}����<�n0hz��ý��+��h�Ɂ��u|�ײ������x������Ѩ����ƚ�iYK�ͫ���]����g*��B(B� ��@&��c��2'u�\����4������ec�b��EOqGM����#w\-��Yl�=���%�m�:t��]	�`�[��B�?����S��S�J�)��ϙq�l�i>ã�i��"(J[�'�y���t�׃`ha���+#�1t��\U���)�*���;�,��Ε�%$���\���q%�G��z8�UB'0�a�(���R0��$h*�(�v����ȹyĶ������{1�p*'���4C�ƧZo���L�~ơ������w�cۖ���p���'�7��LLrњ.�CfF�oiD|�Ь{�Ga"�_��t�+�r�+:~�dק�g?�x�7"6V�:)� ����#Y�͖08`��<V9�'�5��$���֤����o�:Cr_1�!�Z�YG1}b�^��4��|�C���;<�3ۤ�G�� �Ѫ�� �`���kI��q%#4���Y��.c�;@r9��ڍ<�kz��O����p��߶���]P#����Q�͡�Dfs��L���%m�?������_;�<�h�جl�n���l`�-��t�  b��[��t]���!o-ŧ	��=�L� ���<?��!�}�j��o�'(����(���"^�*9#o��/�eH#OjЧz��o�o��3?1��\��Qp��c���6?��oS'�
� s�
@i���4���첁� �λi�4 ��p;��ړ�wx��aK�H@f�N=�'����t�C����B��`��X�l���5X�sq!4��XG�gt��
b]g8�� NJ@=��s���\ǫ`�0��R��^7Xȸ����@�r���`V�dz��b�e���Ih*���n�1&�_��/�\E��W��R��m~���r����_#�B�U��!F��K��������?D��ҿ�A
��+DHa9��c���eg~�L�X�ȧ�-�i�ۙ8��A�����N�X����4��I��޾��E\�P���d�9��P=��DUoM0sW�U���I� �;Z��V|p�	-���3j{��a�8n�D���3�0OO�ː��ؼ�E��i=����?�����#,�_O�i�%���o�~Ն���OpX��0�vs�~U�\��;���V�6���+�׉x�LH}"W+�7
}�eAg��|�_��a+|�J�$�9V��d�%�ږ��@x��f�I@�����D�{pϠ�h���)�S�*q��^�1X,$�3�7I�Ľ_��,K�a�O��D-�i��%�z7�P�t�=(�TT����fEʒ`e�)�������aŧ�r��k���D����Ѝ9�g�C��aޏ/2;Z��������s
-<�JJ��b��*��ߔ�u��N�HR�b
Q k�KD墥���c�ְkg������"�n�i&x*8��/�����=��]��
������m-W.�g�L����K�P��aOp�4��z�jyϴ��9���tF=͸���#Q
@�_�EcG�����./��U�D�!��O}V�uS�r�����H��|����n"�sK3��#���nv�HD(5)(��r
u^��CJ�@���D�	��Uf�cY<��(�eo����L%Aa��􎹲9��Jmtk��U�o��ے&���wi��V�cU}-����w����K�-#r�v�����ڨ`�●��­��|\	�oCn�)Ԩ4�K��k6��.K�?����m�"��;˵�z�{_KzC%���)VAr�N%��R�K�����h~��^%ک;]9�V�j���_�WI�/�[bk%{�9��EV`�;;qL�P��-��`ٍ�0���Y1uUbo�1$�1������9���yI��}����T�իac���8�d�k��Kv�4G�/b5�� J��M֌������>�h(C{ڎ�}S|���fC��]�����[`H�S��Z��T���7��"��܆�ø,�L6�N�gkk��K���Q�R�A���q))Lok��_`�v����qzg�ֆ���kE�hP&v���^�+�:���rd>�>S&{�x���f�s�W*2����4�![�����H��,����5�U��x�~r�����>�J��W������[��g:}��S{I�%����'�R���.2(��^�����rי��πl-�U�Z�i�Q�5����e	�	9Ա$ ���Mx��� Y<���tF��w���X�o�=�X�em��};��$�N��y�ͷ�~>:��Md)
V��p���j���O)��f�Ԩ�I.�G6q� �ݸ� ��L�hd7��^#�=D�m��Գ�����h�/�0�I&��Ū7��sA+4���m�I�؎ݜ������]�WZ�ʦ�}�L :����O��)x���5|@�k6�����I������6��B߷��YF����ěx�V��x���Pon����J���R�f��Q���O��ܛ[��q��X>��9��6���.ݙ���Z^���~T��	B��e��[x�SNbl��ԨW��,��_�Q��S�kʸ�v�/�Zi.E��ܾ��Ё��(�F�{�V�:*NcD�luŤM9r�!2�pZ���P&�T�+ܤ����+���:�p�crf�����9~�Ǚ��6$nײ������3���]�r�bA٫�I5���WL17�0e�l��j3%t�M��4fF���#})wE�x�tݾa}\����|�D���<��I*8���<�jk�j�v�K
)�)|M��o�+����K[����_@�Y?��x(DcW��zK��V��2LjN7h��ϋP�@�r� �����!pP�.s���m�7�"+|	@���&��-���/�f�N��)=+$�F �}��7����gأe���b�Lp�[$,���DdX���I}���1�c�t��*��[�����~|�4s�j��5�3oE�֚pd�3�z�+�&d�ũ�E���W)-�7��]�����7%@tm�-�*N�@����w��������3Z�	ϱ��jQ��Ɯk���h���w�!)������m�׏�tf�g����c	�3��_a�2m(Yg����ع�H$�,��5�t�*|R^�Z���%Y���^�,��=rleKD��mS�P�`H#�F2��X˴'E�,ׅ���!�1�|�t��v`��SC��"��eʖ����6�δ"�_S�g��;=�_M�J�}_�E�^��b*3�� �t-��+����<tp��.*Λ�Ή�ob]�/��k&F��c�)P� 0-��%�E-3�6�>��m�Qkjj5#�n�uLy�[a���)�Y��@il#��}��Wվh�$�
C�v�M:|V����q��Oî��[�O���.�����D�I���8��;h�i[s����`������Gш~�>6��9�*S�Gஃ`۲�V�Zn#�t�h�a�l5*X�/G�B&��X�d���D[	�_m���P<����U���@��l�t���Vy8<�ƚ�V~�r;~��=A�������D�^�Λ�	�/������4-���MW�Ȇ�dtXQ^�ȍ�V�G>~&�e�;h�pn���MB_ԝ�R��]�����3�fiNW�}}X���҂O�y�����L�{$�H� _���+�{MDy�k��ʷ2���!�7�4�X�Z�C��|�vҔ�]"i�E4�}��?l=�V:��:��@��?%�`Nv��[���E�}�*׷�Y^���N�N���xC2LG�+�vD�e.4M���� !��J1�?X4y^F���.'_m��}�=hba8YL�1���3�|��NŰ����'o/:`��(I���f.M�J���'��	?��,�u(�_o�h�j��"������&z�*{��Z�[���
����m����#�ffY���d,}.w?�AJآ�7g�^*�ڿ�]��/�a�Wa+z�����Q�1=&~{��.+���`���M�9t�)e�{s`�� (h#�o��,�Tc�)�EI��� �Oy���������������ֶ�c2��s���ay�'�LP���݇ۚ��G��n��(��N<� TBu�LѰg�Ϫ��rA�.D�ZY��P��ˮn\1[i �#��S�L�\�^�o.<-^ �o�O��	z�齦?�o�$����<����
c3k�����h߁sX~�
yvwO�	�N����U���a~+�[� �������j�T�t�튵|�!���W�/x��l�N�6��3��(��^���u�xd�4������a/}��0����>>yWM��m�d(o�
R�O'8c�b�bC�=�����`��tE�|���ŗ��'$�Q}m������h2�}�0��߉F���jaGC)f�e��!�P�$*��c�%���LQ�?o����`��\��k��)�7C-��o{��ga�Ò�1��ʕ�Egkl��9}�Go���CɌT�hB�_DM/�������*o�@�ۚ����2�"��S
lu�Bi.�{y�t#e!$���%�-|���$���=RcG�k�F��
ΘԮ�,!�n.;h�͐��擿��1�{w��n�%�aR�1���`Ì��D��Σ�Fii^&�	�	�UU��|�1,�t���:��+�eMG���X���)�.����������F?�*N��*{��P��aͶ�u���:����R;S�*'ԧ3�$[�N!?(�����Չ�v��Ǘ��?�﫵��X�Z#;�x��N@��8»�:N�N���Y �j�!Kt�JW׃�Β�=�S�o���z\���WN`t��x\���	?�3G��M>��%gjG7�e��Y����u�|�$�D������u��f�`�X�F��"��tcx�r�;�I%���܆�EM��{���l� �g�;81������\*ٜ
<���5���2��㷊���� �5�0�N�!���_�*��}\���4�J6%��1IG����^t�65N6>���]˼�)�w U�(gxY�X1˫;vQ���Hq�h!���Y��K�<F:��-фu�� 2qv��~[������2��.��@.qmr$30�����mp̈�C���>!�V]��(��mc�X�5��I���ȟ/w��t��zο���p9�}w�^���&���� ����[��fI��	�nʮ'wJ���noM�h�-Up2�zf�]_�	�lc���gd'hW�]>=NO�a��9LZ/�ԁ�����8�Z̃ާ�a����RTڇ\�M/޲��?+�G���a�/���T��F�9q'a���AP1�V��^��,o��~�����ւ�n#�h��r#�pV����H��}w"?P[��yV�]���� 6��iJ�w��UH�������������\&	��;�K����@�j��D� ,��\��c�C��?q� "\�Z`4.s9)��iM����N9��e��,R�����Hwe:���3�ws�KH�S( �hd��|,~��$)4��3���,�����`'��~�1��pV�έWj+dIf;�u�x�,����C�
���:K]N��(�j�����*�����0��z�w[ν�y�d+h#�ol�.ω���l���ؕ%w zIƬ�)�<�lǴ0C���nO�_/|j���v����0�
2��u��^48{���b5cV/ɖs�Wة|�:��m��)��p,�W��X@���|9�˷���m/-s|�5ۗ-�������ك�('�뺏���Ǿm�S�8�&�&�C0V� ���W�ԑ�V�!3��
���������wJ���%W�@l\0�8�hZM�h�6^~�t�c��EΩ���!z�IFr��O��l�"���8��T}c}`�K�Y��L�g�U�]�3X�G�U�.>�����6 �b��-�+�5����NV�:חcg/�3<�4�i���l*���9]fw��d��2�8k`}�l�]�	2������?��������W��ggB!>�K��w�>١Y;�9kװ�
)�= �	Pt�(�m��yʰ4:��(X}g����}��@��YF�)�R���r��:{�X}��o�Y��ؚd{�_��o	���"2�'�����C�h������?�Z MAP���-�����?�D�:t�}�a�.��>!���:�m��+v���yc�x]"��S]yV�9tx?�@����x����;�y�U���a�f%X���*e��)�)Z����d�3X��z�"Gq}�����.��W=�=չv@����a�	=<&��F� ؎�t�/Z��65�!����i8�:T��41F�4������v!|0��o?�[��/:wiEs�CTfv���'/�1n�R�u��2���׻̤'��}���;�ؒdd����w�Ȅm�Ȳ�
�ʉK�W�%j�]_�������E�d�t�]0�?�?wj)v�G@�'�]|�5�q���Vl������~Lp�ך_Sd$���Y��߹�9���3�ٻs����d	��
� �vHa�,$���s�y"���	i����&����+����9���z�#���b���B�9���2��~:�B_˔/����]|<�Dgq)dЬb>AZ��)��b�+���{;X�J]-�jm⮘�b;ILAu[P1���J[ѣv%�zT��[?�ދwE�X����臲�|+.�2
!�J�9_���.l�@�̴��;uq�c�p��<}̱�?�� � x��l�L�9�'�6�$p�}�vϩ}�=��޵�M�l]s����E5�'�˙2���x��-�aU!�l�}hy�%WD[�6�Ì�x��p�VV65���Q
U;c*�]	��)�a��}��1_m�'��T��q�7�^BDJ�ݠ�<'�3�dTk�w��*�M������-X����G���f钤C�ӟ�������60�F?��p������]a���>�fW��է���	Z\1�Ŷ
e(n�n��*�0���)=&X�pJ(���~.�G@���KM��5�� (�p�w�ze��}:�� ��Slq�y�t�4}i�!E�5�"���o�4Dfsk���/ZS���1��{@����~���z9ި�.�|4�UNg)Z���~M�R�<PDZڪh6���H�Lt�����vS�u-_M3��p#7��ƥK�ՏK�~W�8��Qzy���a�.���޻	�������o>Q2$P�K��ԨwH]s��@��˫�<+�"V��?�5��M�ϸ� )����Aij?�V��t�ة��J�چ;J6�zf���}��Z���p	�)�8���F��7m��NY�j?$'64��_��t�(�;��vf�(�dո'�x���n��9��CvmJ�Av�i��q�k���}�����f��YF����7�M��z�o)�.9��H���.��)52�6Q�C2��,�����n��F<y�K��0>�Y��&S��0�fܭID6i���D�=d���wU�'��e�xԚی]w��+΂9)a�=�f,ݍ8C�j�Y��Y]&
v��@���˧t���G=e�a��c���>B������[��'����;�Q]w�MDZT�}�h����*�Ȭ^`1��i�Ɩ�i�D)ް���5�yma���l=.5Lc�l*���6s[+L�S�y�i�	��:y������u�8����C��X�K�.ӱ'�N8w��5����p� ��8F����V�(rk�#�mZ��
-C^ˌ^��	�N���Z�.W�ރ>��WH]��R{���B�|�;�C��%�ק��Mј��C�9�q��[��د�4h�u�2P�ɴe��Z��C���'��6FM���B���H�}p�����b"����b9P�\����n1Xs��RH]����:!��v�P���e��3&%��O�1I/>!�s�9�r?Qș�ʮ����L��Ӎ;���X��a~�H$�[O?��9���.�;��ZKIK����)���mu�a!7꧅DL�`���\�o�DQ$�~��h�-�`��q��̲yK�@	���+;�d�n#�/f�n�ҝ� w�Dd˼a\yi#{LlC��<��CN�b��غb��b%#%�g�&�]��2��?4��m e�w@#wQ��h�S����3'�d��@�-:mk�W#G�F��1�n,����S�W��4Rq��Cf X,�1�(�O�OҜ;`%�GI�^=إ]ԛO��z!b̨j,���)��-�T[�����˷�����S�F�Ͱ��Z@�֟��#I�Z�H�J����|��e�C���c�n�Xͻ���d/ J�6N��ęvަ��x����ޅ��?���H������n���5P:�6�$Մ� Y��IG0�6S�C �d5�7!�K	p��^
��l�W�4ܸ��|a�bj`'S~ �I/5��כ��2�8�g�rǬ���?���5�T]�6��٤A�L��&��n ���|�z�"�������T�_7�N��+�K	7�e�LBQ-�o����2nbp6�徊6XO0ڎ����d��W�Zgz�/�RP������H��Y 0�&Kz��\s��x�O��=�H�KN�γ-a�&'ϑck��N~w�5�ڝ���p��4J��L�a �ര�6t��LE���(�x�%v���X��e9���R�Ҁ~�ymȏ���
M?'SȆ/����7��̾S����q��%uJ#Nd(�_�C�pc�`_��4]�Wp�.U�_u��a%gj[���g���Z[a�ւ��$Y�"VJ�����
�\������լz��kE4�m��RqD	��6�-5:�_)��冢ϭ����(�MC
����]jc]���e��R@�GK����4���)%���B�y�x\ň�q�!�x�H�\�����_lc8���Ë��A��<C�@P�|�E�y�4�r-B@�([L�\�wP�#�5�]�J��"{��,�FEӡ��8�p�KF3����z�ø��S����DGRo��0 Ѝv'W{DI
d_'I__Z��SB�$��w}K�o�%�%�h�
��Q�C)�H�(�����$-'u/-9����k��E�. ���9�|^�Fjk��Y��|��V�Q��e.��p����k{lX���¼�C�>�!�d���ڤ>
�f�[�%)m���N��Ֆ=�֛/�h�Swb܊k�Ԃ�!Br�x�E])Оy�&l[Dn�l3�"j#І��/n�T���Gٰ\�~ƶ�A=`�z�$k��"�L�I)l靖�d�1�� ��cg Eu����h���`�N�+Uc�l@eS3�)N����E�H6}��Cm� �5�B1�A��~�x}��L�~�cks�E��O���H��r�z�,7�[�t+}����v�FL��iӼ��FSNH�C�t4��*��%�ϔC�����W:'���xF_���ܭ�.�3�=ͨ�w ���L& @(�%s���.ϢW�*���bn4?njY�^f�����-�^L���b;�s ��2v�i��!Ͱ�{��\����y��k�6��*}Չ�T��.�ųh�AA������kp�ޔ�p\��U.�N}���|^�)�a	�>��ݺ�s֢��;RQl��g��(FCr��Xp銚;-��OF��Tk�g�R�@iP0}�����h��-�)�ޓ� �5`@S����*���.��:��D���
שbL_O���(��M��ŔT�Ԁ���)}4:�T	���9�VI�ٟ��V��˨�����ņ��NΜ|�J}��f*�j��1�a��P�!�0A#��Ȇ���e�p"
��q�J���3f �)�%����SL��b��ү:P=���?!�q�=�d*�Ԟj�>�G=��T ��v�BB��<���6	-!���.����y��O{�Dp���K$��W�b5��Rx2[�RGH�x�ܦD�3a��V#A�${g�k�H�{�?v؂�y�2�M�ϋK��><>�j%�h��q�Z4���=�$p�$�j���Aϕ&Ȳ���y��z�=�>��^�H�i^��ѳQ��Űʉ��K��f�w1���K(i�P�i/\`�_�����Bk���Ö��e���V��5!ӫ� ��6���c̟�-��o�絃�M���X�?��puF���yy�����ۜ��������LP�S���Dp��T�מ�oxXQ�r�~��T��]����Z���E��o���=����k�N�Ax=��Sԋ�3ā����<��{�@�PQ�E�|���7�X+@V�����C��/-��g#-x�xO�ـ���O~�S߽CE��Ufm0�[W����[�̼V�T9[͠�E!D1k��'e��7���]��YTn�M	�/���L��v�l�BM�ж͕.��?�7�Hڐ�v�1-<=.�W2�ᐡn{nHj15F�6$�~��+�
^lP�R���d\�N���P�h$N�V�u���X� Zt�O4���u$�^�����&�9�hy-�[y<W���j�b
�0��'h>�ٝb:p��z, �c!�,2L9�
��(���:/��n��"M���F�����њ^�?u��UDx��X�p��櫨@�"�H�����u��ω~2�[5�n�&Vk�K�"�!�s./
�&L��8�7Y"E9��:ȿ�c��V�=!��E�k�tO�o��6����A#�/���R��f��L��a&"X���&�m��*9S'�pu`�q"%��L�X��e\�ک��/(K F��*���-�.�/�R
��mS��i�&#Q-�.g�DnU��Y�@/��J;��ω�z��m-�U;w������2��}7Mo�@�d7�h�>#?���i��[����O�&Q�a`9�� жX
g�Mn(:䈻��XAP�����,k��^� ��M���@��ɦx�+8h-T/����d���2l�u��=���Q�Ne���,5�ׁ����Zj�+��g��a����r�`.�{7?v"9��?�xя`����xȾC����
^♰��[ә��jG�^���lkZ��&�=2	�M��S��0Mb�gFl�ݻ�����ץ������*�l#_pD;�w��2} �I������B�3V����q���B� �S��j���d��
�m`�ϟ���F$�q���}݃��⪥�  !��A~�4i�6�<�MԐs�����>���?]�M$�)��݌Xܪ�9#/�	\7�uMaD�9�3 j���g��3Xӄ�)�U^���n�-+�.@g9������$ ţ"n�%sE��k'�wД9����0B�T�ݺr�+g!,`���
�S��S������&-��G��*��" �Ma܍G�WOR]��H���}{��ې��kC��ڊ�Pl��pHD!�/'@�pWR�%���.�\�޴���7���+�D"��)�ϖg�{#. )~��R���n)����ʐ��ġ�Wg�cG�W/W������1QG���� �K+w�M$�
w9���<�t���6���z͂���b�P�~���al^%���)�
�\z�h��¥���RF���3��8U�F���;��Hf�8�RO���ŠJ1�"/[��]�ت&�y���z�� �F*�-��W�@21j9p��*��{ � ͠��QX��"����[�x�N�.��N����; �'ƥ�������>x�0��4��x�xYV���d�@�x���J�~glQ��a����YQ�&��MG|���)��EpΆ��3U�y���&�fz5 ��A����s��C�b:�߿f�hj֚�̄��+�^W~6Zg�Q˷r��k�-�)����Տ� ����Sp���|#Vv�cSEצ��z^�<�/���U�i~6C�J;1��E��,�O�%�rE�M���xv��IH"��w�Ǆ${-@� Y�!�(K��g$�Z�W�B=��R���6L�E�fb{�azp�e;W�.���g���緽��g�l�?�i�_�l0�[��rd��@w.��
�@����B����*V�H���j�^n�R��g�t���9#0��C>��{�=<�<�N)Q�]�X����D��˝} �o������O�o��ǖ�C�h����X����@�DF'�V>�A���m��L>���'�;�b��A�х�ɓ���i���x���E�:.�)^�[���:a��o��ȓ����Q\+���I0'��3Y�t[�*4�}�x�
���(e�s��@ ���r����ԟ�]�
���Z�e�.��07��:�x�M XD����OAd��e��|ҿ�u�Q��q�m�)�.!�t Z\��oF`ڎ��'�ǐ.	�fmi�[Z1��;�`�������伟����MuD5~b�ze�;!�]����wx�5H_��	gn�%��Ɩiqk���'�s�w��Z�H����6�IK�$'�4$:���xP��7�7�?|�IA�B���;��i���l��M�?+47�g+mb��oӡX�	o���c�悇���a��+()�%�=�(�jb�Op�8�|Q�]��M�[H�ӷ{�(�(Eϒ��zp��1�V�����
�U�mj�gFR2���D�����Mw3XJH/b����_U�����N���R`���:H��3;��:�@0��:MkSYM�9�_��}2��n?�H	�)E����5��L��.��_�K�ʝ�k�Bc�l��S	���e3�"��g��E�͏a �&��[y�z	��8�	%P-qq�5�;���(�k�Qc:*���t���gmW+�G����RM��9q˜�)Y�����	��H�F��f��	�J* ���t��!�U��7��o
Hm[ j����1� �"�qD�5�[�|k�!�x��hS{���/:.9.�U�[Y�)'�0���(�+E��8�:��@����o�!�ސ��?��Kc���O�F����A1��$���-U0�T��»<u@�<���|s�q!������~Y�v��8��;p�����ɖ�L� �eZ}���BF���^<�}d'	x@uiZ���N{RU-+zXj<�s�`\9�!G��x,��:�&���!�Uv����2���Q���~@/};N�.���ae��#:Ϛ��Ͽ)�/"�������3-�hփ�й�y:�>�[�"����G���|��Z�����a	�{-��f�]ҟ:�.�9����.w�&G������x����s7�L
�e�u5w8���:u���xu� �b�VV��b��h_d��&Ҋ������k�"4��\�)ݑ� G��J���7I�Sِ-�\��5�jƈ�9��5��/�{���]F�]n���N���!_�|���,A<&x�_�5�2j�8��A"��dN��q��6��۠��} -L�;�3ڪ����'�P�#5��3��Ř֘Zcw�"���N�}Ư�2�oM@�����h�@�ԓ�����cڌ�	C��>N��a��=ŀ���%k�+
��d붉]�^dS�u'�k����f��:,��h�
�
����ӼG��J=��,��_��Ԇ�G��A`�m�ܩ��)y3�����ʦ{K�Fo�C��_P.��C׫n+�!cC�swӿ]⬟�����cq-b����j���|`�'z�D�l�_��p�f��f�J��G�G��]1��In��8�{�n�k�C����.^�`e�,�/[U'�B��?��ɴ������Օp77g�����wА����Fy�ٖԑ(���\n1�q��94�P|0�L��?/k��.I�C�i�1Yʔ��d<�n��gl��v]�:�v�y�0�����Z���b��Z�����ځ7s-��K��_f�;v���IS�"ҝl/����������%�Ⱥ]g>�3!ov�)�m�!�F�%l�?ʢ�R!�� ��CZ���v�����ٌ�W�X*�$7	��>w5&�0�wr��c놋v@
�&��BR	�=�Z��]�g-HHK�jV��ڨ_e�K��Z��ֳO�L=^u�ef:���գrП��R/�I��Y.��G��&|��3�N�J��ϸQy6��Fմ��-��[��䪉(�o�������=_h��9V��۾!8�l!��pz�ѰD��-�^�]�2�-�v�Q5�zi_<bhw��qo2^NFtQX��KJ�uF���*��4_���o��q>9R��u�6�
�hߟ8"��`u̙�����������O3k�y�S�+� �,Pyܘ��|z#�ׯ��c�yZ�ߓ�4�Ȱ��� �P�z2C��y+������H�2��1C�F
��L�6�l��) �ï)�|�2^�]m��W�~���I7�(S�z��@�q"ܕ�
��5By�'6k;D= �Y���D80;�DQ�3�$�ҹ��ŏ��������?��|ZZ�>݋I��<�-��(؄E+�0R����ww�O%���a����s;(�v�\-�(n
C�A!�B�P:�G&Rf�������A䉤�n��B_-��e���q|�t��L'*>F!0΅����5��5��H=���bt����rlv�����s'�X �I�N=lM���d�������Z^2���q^��1�`R���YT%3�(�Zf]ڔ���"_�r^(�f����n��f�=�h�����b���Բ���\j~��Z*��н��Yi�8��G9���o(8���K`��e�Jy[����Z��Pg8��;��K�w�|�@�ıB2p+B����[g��Re��m��`3߾Z��J�'���p�t�gk]M��@��.�}F��{[�[7��9L?����}�@�~�Ӫ�W
�Ǉ���n!�����iO��h��B�y6�H��DeB��:��M�N�����������v�[Au<r�oܻ[[�2
�`��[8��]x��Z�_�,Q�Ō���T���xۍ�(��-[1C߯�I�&�j<��;8 ��ů��˺����IƸ���1�N��iS��t	��%w(�אxR�`�W��Z�CX1�uR�h�f���e�Ma�%�1��h�^;� ���2/pAt��#(;��:�ʠ��������8���W��hGB	鞸�N�F���.�M���|l�C�}��>���-��]�D����^l	)�਀��2Y.������:��m�:#�����l��#1CN�OJ�"��oFE��)¹�!�b1#�#�~8t�s1o�u���D���1+�>9vxn�c�LjWA�[��戎Rt#?lS������6-�H�	��(nq��e�_¦tU������8�	<�t��%6��j��޳��(�aif�]I�QF�`b�,g݅_Qѧ���Ru`��]��z�� �Z��y�^-3�?�=��v?[�r%�Y��|�B�d��O�X��G\�)����Yx��2N"H����f�|��H%�k���\�nݏ
����l2�܃X�OU�Y���k]�x��� 3j�;�&ϸB�S-�#b�%a�f! �ҿ�C�E;�A��:f�q���`���L�y�173��=��3����ZЗ���T����Y&%x��3tұA��m��4@��cf�P� ��_E���T���I�
)%Uꜩ��#.> �Q�N/3g^�.�����9��w� �n[��q�o�5��Z�\���}r�vl���"M��.S�MY���J`��p8����s�
+�PpZ�7LV��$xX�jX��������+�_��|�w���H���:�&UĴ��)�P�Zg��7r�z� [SFs⥫�]cy�x �ϸp��X����i��j?�p�?Bl�!�5&j��Ur-*S�a4^u#T�|�բ�ުf�%z��l��
N���l|DzJ#�e��3T���u�*���g��A-/�i���R#� k/d���� 6Bg�ӔЬ��,[�Bg`�ޒ�8~ko@����-���K�[b>�W\~ �ׯ��^ZIb���7ee�s.m����-P�
]뤪�m���ȇ*����0����X�y�Hqq.Q��� ��ׅ:K*w�|���0�YNu�S����(MRz���*x~��?px��Pѭi����0��Bg���J2j�x�7#1��oW�$UP�_"tw�[�6���.:8�|���7����9#��bZd��F��c�!A�%.��9p�I����/6�u�g����0��U��~ݲ]��J�$���.UL�eF��1�A���3��x����=:[�KN�{�m�L�i&` WJ�H*>�0B�s8}2E{�t��c��~��{��x�ݨ|^��IQ�쑿���C�-�?��E�,k�Jy'l 6����>t��~�6�?�ɘ�#�#���,C~JB���zjG��9�Z��ߚ�hڻ��Q��t�L�V%u6CG�*"��H�x܃��m�iG蟙�ȓ퇕<�H�cMU ��s�˶��_h���˻��­^L��E����B!����Z�k������7��k��'��/3ȳ�	�������Y	|���N)"tZ!|��b���n��CU�����Y��V��!|o~�p�<�$�T��n�/5��J����NA�E��	�Gf<�jd��/�k�<5�L!\�8�/�h]��r6��f/�X�#�O2�Ć�U�qPF�@�V�
�Q6Q�o�z��'�^��%�*n�V�+&��g)݅y�L��JL�ӀS+���I�m��_`�}�u���dk	^F�^kd_a�v���>sͫ���j�ै�=!�-�[,�r���O�u��D���#vT��1�f���[Hv�׋$D[i���Gcg'%D�9�)�\�;K��@�}���')*����ܵz��+B�7�,����(��(�u{��z�\µ)��0(�(eHO��\����G�5A�u)]r �9'n�8�ѷǍN��غ�Ak��T�0�z4Lzx$_pi?	��c��f����"@�K�x��:�t��{�t��������{hU!�"��	`)Ұ욥u�%�˅�#¯:8V%[��kS�Ho56MS�|��\��)�*�=K�ط`_�5�a������X�]�9�g�fI��N�uO�Dq���
��g�a�F�NV �yL\3��X(eJ�7�4�\�Db��*������as�褵��T@�(��gi�W���:Yu��SN2y�G3OO2w(q����ޑ��w�Ŝ!��Dc�N��X�b�ˤs!�;Q �#:M�$� ��$�2���E
m]��B�0+e{q+�����5��9���hC
�J�f
(;��(���OZx`��,�
���Yd�.��!Cf�m�u��r^�ё�!���6V4�8Jײg޳�T���q���Ğ�������p���S�����VZ6��JG�m&m�o����0���0�JY�\�����4�LYú4e ������\�n�Og����	�h��/q�{��zaK��g��!3~� 0� �аf*��XARv:�+�ƴ�JL~���B�&3'k��:w\Pv���62�C��U�V>��R�����sv8��(�HX�J��ܳ&[���3N ��⊻���eO�Q��P�����O�{c葕�ش���V2�ɰ4)����o��G���ӭ��ҎH}���q���\���㖫�'ځ��o,�IW^�7n����J��$[#�!}�GE1�͍�e����:IRA���U�ZY2���[�w���B|��g_m�V.\GC�,�j�[�Sj�\ ����*��6ǵ��&{����;��Ƌ�AH�U�yW���ɨQ9���Ym^�ޟ�O �_��❩G==s9^v�Q -���W���k�cq�"ݎ��z���m�m[B�K"�0�lPS�&7χ�ڹ/D�:�y��A��^pw��є���4Q���d.=�g��R���� kɵ,�^Z��A�O1"�=���럲�|l�u��)��.��%���Hb/��C��Cff��>�\�>i"�!��0���B����<��5�@��1��nr2��b4�$�mU|+�lf��2��K�My����Y=���߰�дX�~���T%�#o�ȓ_!�tF��J,4mSIm��u�8�V���o$ݏ�I���5�� ��re�n)#�;��ځ�CZ��	�/�DKum�%A��Vg�t�jF
J�x2��.Sp��"2l�Z��I� II�V�@f8&���������h_w�}+n�# ��^�	*Q���xn�7:�h���'N+oNW�|PȊaL8T�]\;;�ON S~�NP��{nL�Nv��}�۟*q"�@�]�旵YEoΩk����^2W��Le�-	�ࡏVY�ɑJ��C��e�{�����e�囡��>��rXnD�o1S4�[�n�T��&-����M� �����NT�˿���.�s�W����Ԉ��R���L�$��%:A� � (�CdoC ��C%�&NV�h�Ho
���qA�8�eJci��S����5/\�ث��=�����p' O����G����/��eK9��އ���{�"�I.�	���/�c���2T��$BBm�Ω����vR0�11��=�h�����l����l�?π�����=��1�3d�Q���Rn�-Z�I�{�p��;�=E�-���	5m2���m�l���|�����t/��) �T6*3?%]�������L�B�JT!$fbj^�Me9�\ދ��=�R*~Ɩ��[.cV9��'�mH�?�1�s~M�!y�1���]��a�����d���N��cX�S��*-ꯪ�t=��d�����iA��ǟ+��N�cZoCl�Yy{��2�CK��\�����K���������M����֚B��I)c�Sk�BN&l4O2����Pz!]Ì�HR��=��p����dmj�y��J�ӊ�s6�k�~�3:J-d���Q����mƖLuF�)��;�:�?�xزl2 ݽ�R��ȍ�&�2^�8>�ɩ��n�B��Ïܥ���:��U=�}#O7(�w�y��j��� ���D1���鬈z��hܒ�µ'=�oX����������^\Qa�L����k鵳��l.B��$R�9h~&�HN�^|Ơ9�Š�W��;��������}𿍁큾������=���k�o{̮Ŷ�F���n޸�YnGL-�#���Q��|��y�GR�W����M��G�~!<M�Z��C�ΖګV�� {�x������v[��Ɖ�S����L�9?
�H/8G73ԟ[+�%+�*�P��#��Q�ς�}yE�~`����gu�o��,�7Z}q��Äۂ�>�'�������H�z��<JM3� >�D��EĴ��
��C+ò9���YU����P,6sf�����wE�WZ�2�~4�+_u��S������ځ����+n6�!�C�L�9��C��M����s��q�ͨA��/�2@0�>�,��-m���c���x�pf����F�C����^�9�P�Z�x|�l
�o�]���3���ig����,߼s	���A#�r�\�Yo�U<U[z��C;9�'��wMpq6�Tg��MB��FS��Jv@p�ӱ�f�F�6�����BF��=Mb��l�>J��=��v���v�.�gC掇��R�j=��p��lW��D/��7��B!m��(�#Y|��H`�S%��@	8������uo��.NWv��u��#zǚ>�m�#��☂��w�=Q��"0�p�^�9#f��Ik���I�B⡬�%G;�@"3�;��P5NX}Q맳�,o��\����L�����[tb:`.���\��Fқo�I5[���tгP�,[ì(����m��)��$�]��Ǝ�+��ѕ�y��5���oE)���2�e,(��4�D90�5���0���� �������(�1���l�FK����`��u|ܴ$���>���p��,�D�k��&�XJc#�iƌYx����כ�����炛 ��8v�mxJ��ԫ���w0k�yGh� 5f/�6W0�ԙZ��|���׈Oh�
ͤ�����ަ$T >w���*���_�yS!��oDT溭��鳈}&;T�40�c�,��{Y6 �ߒ�ܮ�Q� d��h�!Y�jC�Fɖ���c#y�XO��\ڋ���k�c&��y�p`�ϞpTD����n�R�)����x�m.9��3&͂�	=^r���r��CA���vP<D�Jz ^�5�:��:��6����]� ��[��.y���&�Ө^pp̤>Q#x�z���H�����]ќ�Fa�����6{R>S`?�����W�8@�kZG�_yʌ0A�Ï���+L���8 Y�Lq�b�yj���y�v����;�������8�c��O�Ji,�4����dw��6t	�G��3���[��O�
u���0�h'��ɧ��1���-��c�	-S+�D���ţ�>� �l2�B�g���o�m�wS��b-?`�����FjK�f�L��c-hu:�/��imh8Ǒ��;F"��6ű��ցy�V��K����㋓�S�B�V%f�L��I;K�w��<sb�WD�L��zK1��m��x8�Q7�>u��^u%0�����`��#�#�U���r3 G7�u�oM�[����5�F���1d^�v��N$N���Toe�Aq?V���#)��@9`u4v�:�I�V�p!�q��ymNf�ܴ��N��������������)�`�ֶ�z�����|G�*:���(����vX�<n�ljp���r 0|�di�p���p`F��W��I�C��>RN4��/���K���pi9�.�)κ�Y�0w�dm7�nX��eM����|�cD;@���\u���CDF��>IS�}Io�S���G�}7����!3u�#�R9���֒�ߪ��r�}lj�UW%}��`����_��3.1,���d�_Fo��ʷ_Z�@�7��e9�\X?!��q�ビ�e��@���R�KN�f��N�{kP��,D�U�.E�-l��Ǵ�Iئ�%�=&�z��c��`s�R
���� w[y��Z�w?��<��KrC�
9۴�C�kl���5
f,"d}�,�?Ւ�t��F��-;�U3=d�V��:R%]�@��c��1���j�Zg��W���uU� H�M�󙑶�)���O\�kH�S����<E˕�ߐ�Ҥ1%A�Y�7���t���&�Dm;��/�MK�V���{Pú���Ǡ.,�}G��t��Tz�C�T%������H*����Ɵ�����w<P�H��'$��q�m���?� 1�1ʔ�;��4|�)Dq�(�z2�����+��`(�e�]��
 2��8�f�#��|�l�j�2�P+&�QS�zR��t�"�gׇ��*L��۵N*�8�����D�|2=��6b�.P�-���l���`�/�_�wv0_�
��wR�U:h����o`�\�8���-_F��L|9��H���۟��kdK(<8b�A���+�{1D$	sk.�W��? #�Q�~��e~��!�,��.<o?�?�>������}8�n'�W
Ya��>G�{����J_�D��pl���K+\�������U�W�j����\�3ˮ��
$u�Ƿ��zk��	��B�����7?�M��^{��ştO
�^?�
̴@���؅�V��={ֵ�'�m���ߴ���ɱ�w���q���t�Z#��X�9.���KĬ���D�k��z��FS���g�/�E!�z��(�w^!��=����|��+u�Ւ&C����=���i!���&�k��׀�����j�_E���$Y;\^D�R�����E���d��+Au�����D�$��8d!:	��L�&uFk<E>[S�t�o*ˁ�4<9@�nrz�f����"CYԨ�UM��T��݄��g����4{\Խ�)_����t�U��&�vU�4շ�#��xA���X_����L`�b��Hk~�0����Р���i��%�R'�k���B#p�Ih���U�?X��3h**�[��pP �{g�o�s�G����͏�
�B�`��W�.���6B�P6o�
��AވF��P�J8o��-��I!ɨ�F�����tm1��{P6�q���I�X��p�q E�@5�)�~�i�(��r��$e+r9 }��u�3�-� �e�c�9�Us���i���.)�K��7a��f'G~���h�ak���p�������v9{�V0��KѮ��
?��G�n�5B��cR#Q�,vqB�}���yw�e�Y���,p�*�"#��`o�� D`�%C��;B2��HT��A������t�ryO��66݁=G�՝�!�э'�(�6$���7� P���)G9����h��L��5��S���4=V5g��P�X�qx:��j��KR':��
g>�ǰ���`��|�{��;�@
���lI�\�S�N��pƯh�`H�,�"8�8,�s�Jy.����իe�Ҟ�����E�)�*�����mc�r�<Ӈ?Ӑ��i�*pV	���q_�\�Zs�W��ľmѐ��[�ڰt�0�������̀	?��3�&8��D�Q������C,lճ�������S��>��?L$4>�/�{�`0�P� Ȥ�KG�Z*Ɉ߽d1�V�h�p=&X*��CX��K�+���T�3C���z,dπ�y��y�=+�d5��~;��ktj�p���Z	�8s�B�\��x����w�hT^L,�v�&��ِ�I�ұ ����St�[
�nn^,�>G����]`vH筀��� p�[D� $��
K,%p�+��FW�cz���c�
�Jhc�`-B�-��[~O��H�[����� yqP_�K�.XIP���81�B�
B�a1��5>�(�(��k�/ws��<|4L�2���C�I�*����?�Qķ��X�ͥF�hߋ샍hp��G��������_+xg�~�B��?�0����N�eS|`���?D^cE�~X�����z�-킜���X�pp�ƽJ�A��g�!7q7O��gΜ��d���s�8Z'�1��>��c
T�ӏ�6>IT���hF�v�y�l�p���?����j���B)����,O��k��E������/[d��R�G�6k�h�8����H���g�����Q��ԋ%��������:Z�W���P�ݸ�x����`�ҥ\�n������ῖ��v�n1��PPLX�����7�Ŗ'ۄ�mg>3���/3 �~kp�h�C�HS
���m��89������U�;:�B}�8N�L��Ͻ�x\͏2��fp��ȭ��>�$tջ���UN�q~��U:ObHZ)�DXL�]4��yw�`�H���l������x�`�\U�w�$Yt�c?�L,㵆�И��#��}R��`G&]jw��o�+0�	/�]7��f�����̝�|;<k̉�0�oU3	 Mv�K�8���&��N�����ڏ!�sG��39� Q�$@�ye��v�{�M���������͉�{��}�����o���0�X�R����V+��f��`s02�@A �������[e�;��#�L�?t"��S:(����K���u,H2HάA4�u?��F�S�Ȩ��\�%�vX84�Tʁ�$��b�?Q����Z$��?������W��m$c�m&�ݤ���tQGN�d��+�'��8K����L���(��厶��5�ח���l����L��0�-�:�X�
���H��C�R�����%z��
�^G��d���cED�L&�G�%�����!�e���)g���s	�a|4TC��b�"�߀�c��Y�a��+�������d�C�E��R�^�8��l��܂��d��}��|c`�FU췺�X�W���xq�RM�t�;2�N��Y䁢d�c��#5�,��~����R�(�6j)��"�߉i�n!ox�$��yI��U� �<(l�����1e�{\ެ�P�8�؇���hza�M���K��͖���i��u�:��?��')s�f*ahA���QB	Pa�"$�v/����Gڭ��b��笛�� e[�z�Y$.��'�^��@GWs��\x)$�G���d^m00f�s�ڎ���M��ѹ�d�eu��T�`@�"�	��-�̉^�0�<aa��-u� �:g��"aI|���V��I�Fz���D���~�թ������E��V򶫔�s�(���r������i���sH��(j�z�F=|��2#.�4_��ֈZ��N���J2I�(h�v���I���=���ü/���KjޅT��h9s3�};���ݳ�5(��y��� ��fl؊�1��/��S�{���񇞮�q&�7v�j�{=�eH��{�`��D�w�ey[u�K+Ɣ��2n����#�e1$�n�=f��Su�oK�s%ǋs��\Y��[n߾c�zZ}],�h�ô3Up����Xf�u�r�Ik���b}���0�'�ݽN�W�̷�7�j�=�� e�n�K���c��$Bw%�P���T����2�(�U,��H�)�����쫎+O�m�;ݶ#�we��}���I>n���w롩9j�d���B4��|C_�4��"��>��<�=�ui�=\��[��#��Y,n������z_O�BN�@,v%�{4@#T;U�|L�Omp0��Eu�m(S����-������?��V�����j�E}G�8�n6�)0b��Lp���u����Hɸb}�ű�ÈD7O���Z�	� ���л�� �q��#Ĵ���:�Ùo:&��,PF8,�lA��(E��%C�m�V�P�ɱ�"�-�����cny�͜Z��;TįP<����} )_D��Ԍ�;�TE�Q�$���CƱ-{���쟞Ti!�[F�����Eg��"�.�,LZ�X�>G\�q��C,6��-����f�Z�\M1C%��!W�Z��g����x����+g��Ei����:�^�̀���o{��j�+ؠ���,�����~��k�I�B����=��g\�k��LU�@M	��	C+̞�LrǇ_�"��/��D����z|�f����� ���2~�u�� �N]���D~���j�-\s��Ԁx:t��_j��+�:�)&	���U�Ҕ�-�|����p��!+U$=��n�(+󋻃�K��vn���51�d�Ś\���ø�]q�C��4����)~����Ke  Fh�DK}�e�������|" ��7��60���0��������M��=q}+qր)�i�����]{_��x�� }è��N�]��h���F��ҹ�J������}���p%,��=k�����p'e��F��Lu��O��9a�x��z��D�� nc�XҼq�(r���$]air_�5J��)h�2qۗ��ӝd��7��Y�<�sog޸����Py1�\��~�D�y�Wh�55�Bt2Ll�q�~���$�%#�7��Q���P]qm�oY��|�v�~�Z}��4���bYEjυ$��u�
�����ʩD[nT#"T���+��կ�es�3|<'� �ux<Y�*���|'s��͓Gu�T���p�Y���(�f3�o�6J��o�e�H�������	V�5^\���iz���S��B1��2��|X����o�Ѫ�ϙ�Dh���ǯ+4zk��S6C/��e`��
~���P��j�P�n�����FYI��%��r�<���:`��}�x|�0��h/�d2�#K��L��^�]�?8i��g?�5�3�P*<8��S!��;��� Ӎ�S��J��*!��>���h�aq�n?��}����KܪG��tp�]%���[I�?��b[-Vhu�k@�><��D���g�f-���-�¡	)� ��yv�k �߅ΰ�ǝ��`�ƶ�JAÌ�f�k.����>-g���^����|]�q��w~K�6�����)��Xȯ����
�W9�>VU�ƙ�43������)�����L��)�� s��פW����@O׷���V����[v�mu#�<��m|B�	��5`7tstɋ��y����Ƕ�=��� g����w*�QE������:JRݮ+5�5	^�6�k�t��{~��o�N����7�`E�?0��#(�))$Li@�a�^#16\.�/���ꁍ��׃�*����c
����ք��߀B������������	��\�Bp��G�J	D�F��c�zqȯ�:���;��t=���?F�uދ�`��>��.�J+"'-+G�6j�M�J�s(�_�Z"3Ȍg�\��	�L���;�}0t�-<~4���\Tz��a�U%�յ�o�� �+���}�O� �d�M�ކw�+i�%.�.�9C8j{���v��R�*�f�<��\��u�4bB���%vP>cV=N�<d�Ӡ�ye��I#��� �W=T�N�yf�%����7	`�ྒ7���e, t�IkCMH�� X�& �ڭX����t���<����c�=��I�E�Ͼܷ�t�Ą,�<`eR=��d>n*d��t�#e�]�gd��mݗ�|�{��$�:�u�YG#�������dE��x`�S���7����6	4���"��u֝��i"ʄ:6�����a��02��^����M�4Vf�)���z�	�AJ�վ�-������n$r�MUA�'׊^�O>�MFl�M��{�L8kPp��Q����@,��8��5���^��)nj�h����~ �H��U�M���ԣ�Ķ&9eO��`�v=#�[�Ȳ5Q��5���e�R�)���_A��I�H�3��,����-;�H!�����M�|W�P�B�L���e���h>�Xȡ�/�#��^*�1if�pp��GY�9W7�:#�rJ����VC�%��C�"uE��F��&@E��܁��M�L1~ �[��a-ĩ�봷0(y1O���?K�SD-�|��D4��#5�������A�N`�!#!��@$�Qn4N��*�������A��D�{R�y_�w)|��y@�q/ީi/(3���&���+�@����qk$^��A�	h�&1�mM��F������8�J����{��$�w�T�tl%�d������^��_AK�-����� Q��!J؃/�#`�3��
\r-��#4�*�r4���~��~�jHk�Aҷ�[_��^�^�Qpd?G��Ro���j����E׈�i#J�%+�;A��Z��%Q5iOL�)-ZFѓvD�U4��&K/XI���7�e�$�%Ƃ����Ʀ�3�w��vܫ�̪=S��'id�䁑W�K`�函�+�wN�5�����
�'/�VK�k�'��AzV+T�oJHn P
�z+����f����^O)��׹��C�xRzAf�R\� Kb��J�f���nBrX-����0���7O���x��q�@��c2Ԗ��^�*p��|Ύ�O�&�/�%�W�!��dR�(��d@Ҩ�
C_bp5�*��X�����"U�MY�1�n3qxZ���#4�>�y���bo~�l�'�Z��w>ɝ�Lh{������n{�YGi�)�k_�̧U'�����$a��x
��{��0�2x6�U�ȳ��r����X�.N��;�Mj	K]�P/cC�U$b'�{kP��&yW@� ���L�6��X৫�}�\�[a��y��sP�2�a��2�[
��gxT"SX�^�K���8�zl�?{X�(#�3�Ф{�^Mܦ�5Pk<� ��8��p�ߟ,���)P����V��ķצ���t�q��ۅ��ߟe���W��M*޵�B��s��������
�!��_�I3��@Gsx"�σ�/3xk
YN�3��Fp��.1C����4;�F�z9��ԉ��i�t\X�<��eJ½"�+�7`��!l+���+�iYA��Xь�틧��u��_�b��b@km�^;��	WX����џ�gV��`��M�3N!���>�#*-�ۖU1V�	�rO-�D-�=�g69^�ʜ/��b�8��4�,	����"��,�H��F�(����ޔ��Ȯe����&m� /��T-!�Ț���Fo&@��_|$�@���J�;��4V�W�n�S_H�vG�!�[���#
���Q�����H�ƶA�]÷�1���o	Z�e�_~?�;ЊA.�OUl�R�
��_� ���|ڻ'����ZeX�/N|Y8� ����7��a��B���j%,���w��o'Z	�,����X�:��YkM���*QYQ,b���?Fx����(��R���K���<��b��h6^��5ݺ2�Hn�W#+�ȁw52[gU)�k]I���D�?� z��4k�5b��J��Qo��ƭ��n��\˛�|0mܐ���ѱ���H�4PHI��8{7��X�$��^R��|�b�F&��Y%�/ƨh�2=��6�һNfNz�FA]��7��:�]���l��ݘ`��o㤵y���!�`��pq§K�P���(?U����ۄ������k�����/����(��y��kk�k�����8���q���W����N|���҅�O�Չ$Qk�^؏m)c=smpvi��)��Fb���sZ6Uj�O9�m߄l��6`:�#4��d~�����Η�
0�ȵ�T�|O
��Q�nt���)w��[F盙W���_�!��~��f5ݻ�+�?��!?�y�z+�	2;��y�]���>��"��.6z�� �.s�Yruo~"]ߟ�t-댃."�Ż�+=l7���n?*����8ˌ��ʲOKW��d��G�(�9�.)i�|����Z@��<�dN}G;ݙ�'�N�✔\k��5�oR�+��cV�c�$Zu�J���`�9Hc��f�b����@ ��M�3��6� b`y��<�by�^�*!��'E���*o���CBB�[���S�-�7pp�6<}f`�Q�P��z:a;'�B�1��)'#߿�~�$)kJ���~E$TM#󭣑BM4-�Α��i���FO\�E9�Mbg%�I��JR ����y�	7��]��9�ޤk"��|��4Zz?[���ߗ�ՋÂ7ݛg,;vDo&���L��G���Y%��b�e�^�$]���\���i;�c	C�>$��Ԭ��q����4\�D�Ю(>�˽3��V#�U#w�Jk/������94!��=M�j@�%���\�Mi�8���	�<�r��l����QL������K�J��Jӧ@\�gO��R�h�cR��Ѐ�D<܊�R�4O3\�܎%���P�$j�F�寓 ��\\�I�8���s���V�썜��>��c#�ك��L��� 
)ݓ�}4>�mF���d������M�\���F��Q4�1ԃ�ulx��(�0�����N���"�PN�ٛ�J<��gnP���Bk&�,���X�?!���i3�%��wu�%'�e"����3�+�_����c!|�Hԑ��A,����
��@�6N��2V��d�!J�����"F2I�V���~��~>�"4?z m�Y�A����x�R�W��=��*��aih�9RȪ�.81��aW�nZz�^��pͲ��N
\���F)#�q�}ZW(��\�:�w�՗�MN��3��/G�Ph����mIh�W����&pײ�����
����wd%/�(e$N�;�$�tEܮ�v8y5��T��v�8��33d�?��퐉
�XMw����l�&qɁ���V������.\Q5��	�@����ouID���	�P���Y.�u�K�UjKe�^�=�]�&�N.�>�1%/�.�\S`�v�m�*N�d�	�D�Y��o�Ǐ ��S��(ҫ�b�Q�Z�Ǐ-���d��!�z� �q*>L�u���8����{��fL�A}^W��6�}#��3�%)���p�a3V��k1%(��yv>�'71O�'2��	�m.�DK�ý.a�^�ߑ��O�K�` ����m���̻̈��e�8�t����o��;Ze@�у�/�A7�]7gF���~���=>M���@]��Tx}�)�ݠ��{9�o�j���F�}B�٢��d:�ŋߋCB� 1n��ZU�3�g�9�ָ�eOD?S9�4K.�'�=���D��/��z3�ؒ�V���z�ە�h�'dW̞�}UW����+�*��6lMs��,9	�ak����ڲCGŎ\�4�ѭ�(O��@q2D�u2��J�B�Y�?)	���������y�����1�ΛH4n;���>����%�S�0�P�kp��@ޒF{m�2ƭv,�$�r1���O��:��D�#�!I���$A����]�շ}�U��������t�̣�E'8&ߎ�ALņb��-b�^�d=�WY�XT�d!�mjW|���hr�*��.v��Ίa��{ry}�qF���*>I a��Z�}������#���A]T��_u%U�� �?O<�^���< -���U#�l�g 4�N���0n���,����Ci������[��J|�hDmAQTK�lÄ4lH1�1	��PX'p����/!�,�u�p�]��K���4��2σr�i>��Ev�>�s"�,��T��QBg��/S���d�P��,'}���b��={�/�*WF\.u ,Y-Z~�|m��`ǂ\O���%�|��M�	�]���fDtc�?g�a$T^Ѽ��W�ަI�6�K6�*4qX�&�L��\��2KlU�Ej#�i5e��c�X�E Ýۢz~R,R���lE����/9�����58�B�>�˿ j�K���Mz�?+qh�Dr�g
�<e�ŚS���H� ��xlV�:i���r(b���)���bG6k���n� ��QO9faX��O9z�ᶑ��WE �_Y0�e�/y�3�]"�3��^iwY�[Q�ݑ�����p#���"��ء��N7Xb�������ϑ�$g8�԰m��ڋbɜ�;��%�h7ӽ1�Ԉ��u@�9��SW�� �:�6�z�5?�.�����H��2i�Nj��V��q��p7�`��k����mq���3X��1gk�s־u"�6��oi�`xʼKxW����uP�Y��O���0��g���Sk��Ki���y`��
�Wm��<M����[&��nȺ�R�iYS �����Vn���;sd?�����[0.���PW�rxpw�Wrʢ�`&W��{�A��}�VƬ���~M�nS�1i�}l�wh�O^ش�wbr�F�{C)a�E�vx|���,���PYE�kg{��7] >��'E23�E�nʻk�/�jCNo�y�$��К�^sS��S�Т|0��]#����$K(6��'h�=�t$��܀%sܶ~!2����S#�G�3/`���
���=V��m�|��1�Ė�⏞z#L�	�l 궧����4��Z?3��Z�CL+�I1�?����K���(��]��:eP�=r�!��G�Sh��렳��~w��e���j~B�]��P&��C(�/(C��z30�R(������06�!(o���&��=��T��:I8r�l:���^�C��ч�d
�����J1z�:�m�W�����L��QX�uGh3��x���L2_����Q�#b�%��%�\��4%T�/E �=Gǋ�O	lB{�Q	S%G۵�%v�p��B�E1�vjYؤ`���xS-Z�?\�<����@�������+҉s u��3���}Kt�p�B�j�*z�A2�1�zϛcK�+���\&������KL��e�v��4ڢSk}�,��=r���$xaR�}��N�ǀ��3�B�#��.�ñT*�#�3��qa�`�o�i��`�O>��C�ᆫ^�T��(�-d�����rw�-��:�a�����)u�%�$˽*����3����4l�:Q-{q�>$j�p���Qt��f[B���-��0��j	YnD��6D��P�.������䃿~=��Q��s�j���u�=����q2/�&���@�����@����΅1Bò��LhXߢö���haX�D�9����FM@9#�����R�LH��LJ�XR
6PRABa�co�5�7�p_x��ŋG�"��ͬ>��W�R����"d"���DOy��9�2�X���+5�4�O�Ҟ�P��c2葵9��/A1N\$���R�B%�ߖ�^a�5�R���ĎQg��P� ��T	@?��d2��#�$;Q��@�ÅE�%����ݝ���J���l�L�u����
�M�KwTe����9�jO����mNJ�#��T=h�Li)f�V�Ɔ "A�7�$I����IQV�+��0��ݕ�yvܾꥦq\>��Y�"ϩ�� ��
v�&Cq�,(2c�p������w��$�!F��o0�A=�A���vO�B{{��!��Ӻ0�e�P�(Xt��4v�-@H�_7����,��gܠ��	zrSŵ��T%a��� �����r)_(Qa�U ��L'�T�(�\���Q��ːV��nMw�]��x�ޮ� ϗgمN� ��!�~�7TPg���`�<w������Ѐ_��(���e��"�Rs5|Dw�*�ǒXH!��*�l��u���q n�%�_<荅�K@�U�f�f`��YC��}�cO�p?v,��I�8�3pE���+�h�%�n4��md�Λb��r�ScܥX:���d:}FlKV$���j�z�㖧4�\�*�U��a�;��8$��b����oSB�1I�����6�c�`>�n��E��6�P�TCJe�t��T���xb3P�����DLe�p��[��"�k%kc�n���s�t�i���@�Au��փ=��M�	�Xx-b�a߉���tx�U��kz)��p����68��Xi�K|�7ﷱиP���AC�b��Ex��Ec��V)_���^��|2/��Iߙ�e5@�Fw�
�Mg��W�V�!8|�����m���Z���%���¤�i���*]Z� "kڪ}����0�5�D�C��^@�pS�^,i��	j��B��{Mr8=w��ԓh'�c|��1{C��ө��v�H�*�R0YQ��3�͗G�m�������<��iS�}d�Y��l&���f	B�`�zd�(�;��-�:�$�jf�/��i� b;���*h�<�5���9���(�L�J��fa�4���(�N�0�hґ�9���Ui񅕷{��� �K��}wp���x�Ѥ>j+���yV,����e��a�9P)����V}T�hH��?@�7��b_c����n����n��'�J��5O�{�i���R������f��|_���x{�����2�w�m4�:[+n��9��A�p]�H4X`�~~��I�~y�rH�֊")b�;�4���A�2L�l��܉*Z����!�tU�j^���+̚���L�����$S�TO*&�z(㯋�x ����nS@��k���ɸ�MlSJAk��[@��(^�'ߜ�����<3����LZ�ȋ����ޭ �o��Q��� �`�K��j�GzwO~
r}^�4P#	��&�QU?��!1�8R�c	�D�)i�"G��G�=�ﻓ��s'���ee���!�і7an����X9��7�W융�3��Mhp�N�B-!�R��q73�h7J��a@�nVo��J���д%��*�m>&���ëv�=��dui#UG��<&E����o�3ϥW�lu>������F������(c�*���y�N�&��*�7���N�\�1�&�b4�[�\e�
��Y~�t%Z��� ]�b)�(+=Kއ�h���^M���G#@�����o�%�#��h�}J�`d&�D�vf��R3�>>֐Xk�-��2@5b�����յ���?U��NxЗL��̭���O�I<ʠ&C�hQ�+�*�5H��Z��]~��hڴ�� �RnP�:��6�4D����s�j�w�Pj����Ue:.��P�Dn���9��{�-�
/?5��_b���nX&"m��˕ɧ�� b�9�Jm�ﺋ���Aed����4�a�FzI�����b���bǖVFX��)�=k޴�cŵ�Q�9/�� �'}(e脍��K��G*��N�5���(��OET84_�8w:��g�ǌ.���aw2���/��fJ��ֱ�����mnc�J���*�-��Ά<iY�mT
F���4)d�����Ȍ+�ծX⾇��j/��ׁ��UgD��ש!S��ݔ��~����R��KA�oK[��C�}@�-8O�L�b�Tɾ����7"�2]������h���FP.E0z �T�H����
�hl��*����Sd�2�#��&o�#v=q҅"U�\�>1�&QG�%!����T@e�fE#{����E.��\���;^I&c'FA�rm6f��Œ-�8�����v�)_C��F����ל�ՒhaH��F������|� !	�I��$�?�[�2^��3�MycM����i�B1�IMDǬ��Y��E|j��c��/��`��ջ<�-��=[���\��/��J��[>vb��?�VI�.�Л�*JV�RQ���u%��I1v�t�rr��e���<+F}��Q�4�B�x��9��U	?�p)޺�Q���z��bXR�;�1�ƿ+�o{i;?�{��}f���jI���{��a��q^=Yz�c��������#�dV��7 �Tx=d&��	�?�U̄�C{�7�`.����U�%~����a֊앫��z粷º"��`�7|�9��CƦA~��&I8Ye��B���C�Z߹6}�*^{������>h�D�t��(�f��Ҙ��) ��Xi��_)`6~䢜�L;��)�����r��ɯV�m'`�pb�YA΂��5U+�1��z-��+�>e0CB$�l߿IU5FZ�y���ew��$]n��?�ٖA9��K(�?�N����1�1����8*�J-Ȋ�e��nT	��Z�a�]���pD�U�>y0!���Qᚪ��ù�|ta��*�ͷ��ȅ��5�n�!�����nY0D������d�:�{F{�W��0"�_e�{��
>R,(��*&M^1,iMJ��;�U��I�.�`����G1|s_�,S���,��mc����$���t�/�}�IZW}UM�Glݩ����P�������ܬ�d�͆!%?Յ�z��|��n@��^X��{S��@�$ҙ�=?+N>�d���;����!,�P$d8��ز�{&�mG̴]	�<����4dV���PM��ː��K��
(�_�h<Dj���f��`�f�b��@H#��88k��"���@T5��>�{���K�5���1���M��=<���)��Ȫ`hh��֊�ۏ�˃�~4��Z�u/q��Y�ߎ{���'U�J!�"Ǉ���|�#񵌿`��*w�!Z��ڣ���&�)��P�8���j�Npa�+�Q�?�'���d�b*m����J�ldd�XG��w���G+��}��j�i>��&?&�	�^�m���aB@,\PV9��"�?q�u~@ﶂX��~n����:x�8y)ؔ	��L�Vֽ��ԉ0��?��L"Õ>��a�p�ɜ����_=T!r��A�Bٰ<��3h��`#��,��8����/l�F�h��!?aN��8�i�[�\mi�6Ϋ)q諦+�2 �Y�pr�n��:�n��%���:C;Կ�<�5!9rU� �ֈ�)>�����!@fSwfiCi�y,%���_E����|�Fh�<�8�����Ogψ<L`���fZ����z%i�-�
�(��H���4���g/�˼��K-[�j�ӱ،P=
$��-\^��m=`oYU~�A3	pR���� ��<ƿ�_F�q�q����-��Ԟ\I�A��CS��̏��4�^���5[x\~�w@բ\���p-ө��hѲ��=�������2���|U�<n^U�����(��+ũ�8ck��z��� ,6����-��~��Nr#WQy��D�4���&Q�>F �����K��S����sy��
��d�S�-tV�z3f���!zU��R���i;Y�g��1\��`��[�坝R�Æ���ȡ��{M%�s���x�87)�ϕ�����u���Y_f��5�Z�6C����.�-�<"JGE�m�p���ϭCu���X���w�LJ&���i�lWW[[8=:�X��f�`۠��$�o2DP���WR��W�8xj��1b�Q��ۻv�����fSd ^Ju�v|��������lDŝp�*s!����No��x�F�T)�d���)V�bP��e�����0	�-}u�>I]�ò ,/��Mupڲ��hk�ۢNm{R�N��*O�O�p�������(c��a~x[c��-~�3�l�z`k�-����L��"�{��p,"T��Y�S���p+��J���-l��'B(�p;'=Ejg[���:u6���%��l�Ԍ��GQ`G�T��2W.#�����+U�{���Ō�w���2�9Dwe���0��PE�=���4�KJ���\ܦp�P�C+�qc����
������A����O��=����jn֔M&��6e�X���7�IW5�x�kx3��Y�����F`��+ϡ�c-�����b�;"�Ƈ��R�	�&�����
�%k:P ����\�q�fP�ѯ/��-���: �'-����{�$�(n�hT��Z�G�Q0�=�x��Gq+O��޸����>�����=�1�)��!�.�;�0���7ي(r�E�%�S�Ë�W��Kv�ZR�r�`�c�A�u@�^`&>�﫮��
g���܁[��/�+� �^�'XQd9�awK�tj��ݭ��(����+}�4׭�<�ei��`@~��g����6�beXrv��0�Bu���z�B�!(�p#uQk}���t���sm�D��ʡ7[�����qw2�㹛v!1�p#;%���[)��k�7#?�k�3�Qe�J�:ó���c�)1DB��A�q�K4h�"�>䶤���>�Yn�4	��=LӧRB�#x�˱� ������WJ�r��H6�b��@�%9/js�<�ć}�6g9��B^]p]M���Lc��z�ך�5ƨ*PhR+(6�	�3�ޫ"�/)0��V��<�Mܘ�����3p��`;��I�Pt���{�`a�j���-2^ɷgו�I�'�Zf��i4��IǪ���Ә ����}�1a6p�n����9�E S	|�8�K��d�ʶ�D�8�9���B,�B��pm�Y(DjBu�������N� C�R�rw�L����-A�*��v��Mi�EK�!��WL�`�3}���*s�=���e���v���L}PƝ�?h��y*��q�ٌ�����}�!�)�|ڥ��˞��䳷!���/��#.�Ɉy���@�-%�m��Y3�S��z4*��e�����eϷk?,�#++i3q�ͣSI��<�p
��Me)���t#w����2%���2�F�C��f*oד�SWl0L0�[��P�1�@*G��Q��R`��{^~NQ�GЈRa��Y�������1 Y�s��p�_�fo��zJ�����/�)x Ѻ�����n0h��n�y@�Tu��Q0'F��9�#���v����mݴ�1�\�����-H\���T���9�T��Ñ�YC0���3�ˋ;X3! ��I��eL��Gkx���x�熺K)������v��觵<㷵�/6�Mɕq�7	���S�/�r���`�`���*�nΡ���;7��]������~������1$7��F��[W}6=|" ��+~4��!�4+��Fv��� C�b$���[f���J(
���߱/�i�0P�J�Il4�LB��[���U����ŭ��m�Ė|-Fz!g� ����-.z�#G��I�ӭ*A���8��|��#��ɗ��i��cI]}��v�D�(D;��a�m2j6�p$������F`�m��bc��(X˷�wxs�Րا�E5�{|����ă��~g�
�r.�|�5PR���B�"̐u}����A-���5��F9r���*���#��ةm�P�uE�B��Hy�&�i]ps�a.�	Z!<�b���P�I��C?�aˊs�ܧ��`������6@1�I2q��&���{�������bơ/ʯy������ص?�cBYv6K�f�hQ��P��	Q�@��#��(�DE4I����=��X8�bT�LH�H�ש��x��M���`Y�*
��m���2k4xý4$���a���N�^"�h�	�u���6Qz��=��|:�.�곑����j���F��5�l��˫ۧ�~�T8���n��l1�{.dL0\�����Hx��*�v��ُ��d'㔌�{��ʤX\p�.�5��bi�|��)����n������#�J�8�|��w�l�	���s�Vv��������M�\l������U:��'�5���Kpr������W�氓�����gs��>&nZ�I�7��l%�F��ݜ~]��v���H�	��`�@�P��<�j筨P}��9���\��#�R@u�[�1=I��|�-���N��t�{`)G���_Ƹ)��,�3�� ��Q��ޏҼX%	0�B�>� ����0���e��U�:!���[���Ht_���W��T���� p�rS�?��ML���j��X�U�B'��#G�vL��]���!"���
��m�Q(��EM�24��p�A�-Lx�R�d�YL�;4���KM���������<ܠO{��'�g>���󙿒&�/L�VF���>�,��[q�?8�!BL��;ni/�����}Vd��:��
/9ޫK����g�K��dxRL|��+;Y
&,�M6���rE`P�E��v�з��LX��/ڥ�7�ꍅ�cZ��n~'�6s���������4D��F͹��H�]Q鍊���/�������\��2^�2݊yj�es�ꅆ�L�����f2���p�\���3v�����'?�����*�79B�7�:�&&�{f)h!��c "5V%���%��#��W��!Y�M�Sf�@����	|���f�)��^c-f���1�N��$$Ư��Q�@�q�툙��x{l�����p�֠ᘏ�㻡"�`��ߎQ�����Wx�V�X]��T8��
� �mF�XG]i����I8ib���i:+��rV�C��7Y�� h�X�JE����[�����jy񓾧 5�r�%�<�|����,�_;�, ݼҵF�3�S�/R��~I>���ws��8�b��/��ۯ"O��X$ٷ����1����?��_n腀[0����7��i�j/�ˌ��N�:���}G�L�.�ⱌ����b��=��?R#m�Z^�sC��r���#JU!>�G ���z�?��0Z\��� �aU>�/3	�����b7`M��bp����y�]�e��h{���O��$�ۣ��G��ilRg�Yr$jz��c�<d{p��̓�rT�M&��� ŗ
Qw�2w6�E:I�re�u& ��r�*Z>EE&�-������R���ޓGo�>#��Y������σ=�a�2�����D����D�߹��^S��6yb�H�a��vI�2=�=������d�aS�3s��^~��٘L����m���(])�=L�ۚE��+��YFhS3+_���N��2؅���2��C�D09c:��j6u�n��_t�r؅��!��7G�*H�J�����CZt��s8�W('n�콴���c����G�A�u��������i	�"\䶦�d��Il��0����LxIO��	�ؙ��S�#��m.3*f�p��'���$�Qу�V��	�O.�&�L4*�՞�HoG�~Ϩ/��$&��ι����L������9E� 2����!�z��ˍr���ULE�(�8F��!_���%1�+@꼗��o@i����5Hn�-ދI��XGp,��"���6��:0T,�*����p���ACr^�
a~�����2Si.|��H���;Q�\ao Ȯ��5:��:ȮB���F2*�_��C�P�]�+@4��6(E0�8���h�\�R&<w�*��T��G9�r��3���0U��Qt�����{��߸���Gv���I�<ޭ�ɇ]�U�ϸɴ�ś���}m�ԝ�o�-)G�nk	D�trb[�Z/�`���B%��VP	|�Q�f�i��U���+����n?g�H��m� <�K�0��Q�E-���* (����Vr*s<4y��4D�{����8f���s1@MG�|�>��s�N#�@�^�� �| I�<i'۴��i����Z��ӽ	�4��� �i��&)�˂���=��o@¸ɼ�_a_t��#����u�<o١<1�g+�Ҙ݆��:S[ZO'��R�����:��V5R��Y�@Sz�m=� ��bRK�7��.�yj�G�a�N��a�qq�j�٣Gt�ܯ!�1���(v���gcܹ�����h��E]�@(�� ��j�B���>l��FT�0�5X� ����u��Y�3kP�n��$��S�}��O�����5��O�#[��hNwb3)���ۙ����`�H+���?1I��+e�/���س��I��##3��U�h����}�I��È�|��j/��݈�|��z�?��*�����R�.�Ҵv,Ќi�)K����`RIW�6��O�����;"���b#T7J���w���b����5*Mu(�-��5�-Ǆ�m$�)�P�S�J&U�C�0t	eL�Ǖ�k.;F����cK��"��9EE������L��	�]�Ƃ�a�����M2��;�ּ�:Va%�Y�����v7x9�.]�����+�@v���e]�� �z�Qc���w'Yԝw��]�1k"ߓ��M2�p�~��3ɛ8~��1ˏs�WL�O�݌���	��.Q�֮E�N�ꋜIw�.���ז�CD7IJV�1EJb���5�K�K�`9e��J*�9N�����
���7�Ni%��MU
�H/V�Q�)�.$������� �3��� ��s:$�ȕ\��<��9�z�=}�q5���Z}��1;>�u&��@E�r1f�tU�o�ջ�C��ɍ�/Dn�i�F.��D����fmQ��۸���lS�u����PYJ�xЉ@Z)OT����Icr+ȟ��7L��VG��$�a;�L/���D�m��B���^�PR[�����q ����W�|Xy���D�+��a.�c����h}odp�H���,�^|4-�:tI�2y�Lצ�b�=�~��G3Pe��~ZW��/�'��O`����`���Q'���\���n��>��|�9��_�s�hZ���	���s��I��W��+���5+�IU��-�PƘ��HXjd�Лm�r^VƇl��"g �;�Bah����,�Y-���&�!-��<����F^�ιN��]飆�	7'(�.-x57����1�%e*�p�]S[䵡G��L��(qp��e��\�� ~����c--J:i�t-��ZHC\��h]YWO*����k�y>�EU`'�h�μ@���� ?|�A�Ȼ���"zD;J�.��2���P�?CR�FX���8~� `5x�ǀ�Z �	!s�z��M��
��q��D�4|%�%�a�&��?͒5�](H�7���7�K��e���cń�K�A��T���c�p�˶0�(?gi��q��jɐ�-��j���cO˨�\1�u�w�9�6('l��TP|j;z0�6c!���EA_RHj]j��gƖL�s�Y��/��_H�oX/�b7�����p�@��.�5@_[���YK��氅��C�J�"z���I��%v�w���Ɩc�QmV2bC���
�=`����Kh3~W_����ZJ(d����R�+��p�s��c��B�s9
2�\.QJ��0�KC�+s�kz�z�}����E�Z9hY�;ы&\�.�l�kݷm�#�H�<���>f؀���%45f����(j�F��Mmr��K��#\5������*+#�j���F������Î���5��_��o�O���
��� �9)�;�?��-gs7�O~�Q�i�
��(�-df�A�^u�����\�;��D�<A�d�ۗ����B�:�"��z�"I)¸&�2�1D��#��tM�t�ڃ�\6���W{�_m\M�G�_��EJ�iݎ�ʧ�7pH����oT �zSO�
���Y����6�)�!i���R	��/:����W4�M�0\y�˫uMZ�:�e�j��}j��5�bj�]j
,aRh�t �e�/�J�Zm?'��	����뵴
�a�X]t�u�^ԫ (���F�i�3=	�	�F�8�;|�@a�c��1�G{<�@��N<p�)j6�ws0���R�"ES����K��p�����>>^�vKa0�RՒ@Vru3�7L�y�?��_� ��H�0�9��U ��9�]����/J��"y����we��DΊ�c��\��[��T��iy�Fe��.��qx����K�f������rӊ��[���"��>���h�k63t}U����9.�A�
0V��x�^+��O�����:+
'@^T��X�+�Xz���+�mӷ�M9��a������*��<[Ϸ���3��C6")��6u������r�ѐ��J ��,C����p�I/��ސ���I��!������$����QM�o���s�r�<��^��}+���Ԋ�A�&���q5�t�*T�,
&X5X��Гx���R��C����R�����(vts��^[!5�^JPVA�����  �Ȭ���4U�cpdM�ˊ�XN������P��tp&��rD����\,��*\h�{��2�_%�+*��r��)��0|�P�Ir�Rr�7��{mF?�"}���׿��;&��bN��L�x�b�1;b�#��#����M[p6�I��-$��A"�`u�T��j4g(R)��Ȧ��%�G��q���[�D��<1س�)O��2<�2�c��[��${�Y�U7���%��{ߠ�oT�J�|�@���>��aJp�`�vVA]N�c�V��Rh�Oo�xz�8Ԏ��1��?Ϯu��2`�a���H�
�Ҷ�X���J	�ط��#��ڙ��0���\�}���\�8��5X[3�#�
z:Ɛ���V����܇e��卸���7|H}�`w\t�S䞑<�8� ��4w>t� �]We0�&F��(I���xzla�B���1|�
�B�G�1��/
�Q��:�Y�7�+:�y�e��� �B�/�c4Y8��bS���4����9>a�]!�-���z����L6߲�!h�C���]��I�8]�A YNg���M.��x��VO�O.�XE\�b�1�ag�s��܄���A0K�z�@ĝ��#�W������4�&v|9n Co����ul_%�,�;M�i��V_G<�ᇄ�K����y�>o���.B1�O�n��T���5mN?�o3,5�x�!h�څ[���jUq$&�o��`Ly�}�񙈍֧'R���v*3�5�6y���'���*^,^b�$����(�~㘋�=�hm��4F�panee�]ܝ;2.�/?j'ݻ~�
;$������~l.���@X�F�6 ��C�UJC�j�aZ���V�6�K�,��K���L��.*C��1B;��1h�!�ǅC,��&�V��L`�I�M�����Fы�K�-!�'�,N��gJ��|���|��CԻ7�n��z��\U����n�&�t��i���"�i�u��i9���@��Dz���7}l��_Je�8�U8���'c�ƣ�1�Y�f�oN�z|&��)��y�������sb��n���4�-c
��Iw��'[��<:�'U=v���j�����u�w�u��̅b*�D�Jh��ti�
�!�!Q����} �<�(l�}�}�;}{��V��Ӡ��C�<�L���"��)м= 5VcC&6��0�4�Ӓ�s�*�b��ص���NW�#�n�"���|�Ce���#ca����`U^!aL#X��萔�������;��"��`�ո�؁����Y�M ���ߡR(�$�0.�ޥ�g��Y)I�q�sd>�G0u?����u@N�e���:�p��` X��\ѣ�ҵ�O�����"�_����%�COQݣ�;Juk*��Y�K��mV��*��D�u4��2��;K�rXu�eTT;6����:��yΏ9eT�.�<ҳUm����i�s&q�2s-�@pY���o�Aɫ�!_�>���N��
6"�i�^�^v`��
��/��BdE�K��s��zG�F4�s
���P��4X		���V�3��P)��f�<�<�hD�5��rёD��M<	�������Afh�r�s��%�xЅ7�9	�6oMqv����8�3�G��	�Y����R
�;���h��Iٞ>O]�W���i��y)o��,�Wg�t��eWwWʬ��|��T�������}!���Q�)~d�z0Fr�Ph$%Y��\gr�N�"�7{O9�g
�ѵ��T�]m�"
�B>B C}h���g>~�=���B�L��dv:�vT�:�e��-��u�D׵��H?���@P"�7Rm{�㩅�?l5�;������8�'�0:&BV�kg!���E�x~,��t5hE1���8�D'1\E�S�����3i��!v��S.Ú*���m4	�z#n�a~j�b;�6:Et�'�)�$֛���S�H�ȷl�Arᄊ�mly�����>{NZ��c`/�ܶ]3h2�l�q�����CP��k%yq�:�C�B�$Ed[��!~�?9l"ȇ(/]�p�	GK%͈z��������S�u;$J��@����B�
-�����a^�T-v�"\Dad��H��E�?��	%�@��V�E�%����a����ݘ;'���d�]~��+�8W����­�r7�3�H��2*y�%V���N��p��df�]��9\�s�p䠹"Cu5�=
���(%Hi�"�����h`x��I;��BA
T^��}R�\ci950��;38*��!6}ЗsZ���)�nj��������;�^v������?�K��B�Ú<dK�V �7 �ʲ��(��I�����^h��L�=���CD��a�Sf��N�'��X�1���	��ې�sp���R4�������[h'>5��;�'LS�YB�G�~q1w�Jc@a�Lo�_�Ij�x0���`F�gM�d�-�^�-讬5^;=���5� �9&�z�s��_O�Of	 Q�q��:�g��H��fU�H+����g�V��+�X��pù�i��E-�
^����L�+�j,�f�V0�52T�}U�LA3ߘ��u���j�l�����F�j�5�$G��jq����/���k
`�d�0�ZH8O���F4@-��b��/;��+�x�W�����gΕ�r���I(:*�1hU�t�6r��Ɖ�ԁBw���>T��k<\ v����k)�� �D�'C�.W>�ao�jo���M4r�q������k��g9��*�M�X�+����A������=�&����8v�i<�I���ȡ*f��2��1��&~SC�1jv��oYy���D+����lk��J}�6�e[�ݚbs�̜#'�ϲ�G[����J��!��˧�:{P�%�v��qS,2�jL����;��2��0;�����;��)��(X�zeBc���T�!���JF�N�
Ŕ����e/�}���m6۸�3�M[Ky���$F ��R���pa��7n�qc5�a��v��� �9�T�"I�8��0�/B]&��9���p���ʰ\� �E�E|x	`+U�|�%�1�8����V�_�_@wir�Y�*��gL�#��O�����Vh�0�ev%�k�� %M�>�����c�>X�ʍ3�%�=��1�[�@XЛq7�D�t�<�ĉ�3F��'��dS�i����"V<q/���e!�RKỲ]|��l`����1Q�|�Im�>!�74��~�?0FG]�>�VNl.��R�A]F|&K��]5T�b�ɗ��ǅ��k�0A��-v�)q۸=hP�â40�+t��є������|�y�'V_`H������,#ؗ�T��Ơ.��Y$�d2/#UC�)�eN�d�>�&i��m=˷�5�g���2
�|����Y�t@�z���ְ�ʦ��- ��=�*��+���jӪ[���C(���l
h�̖Ƕ(u�"��� ��_�}C���4�m&�>�_�!��}�\���f�s��)qai�;mO·���{ ɳ�A^�̉1�m�/�a�J@�w�^~,R?&�	�6�1i��J��)��9Y�e$ϔ�� �`�����t6�k��16SL*�7|��a~.�0!����)�p�ɂ~�q.���e�L6���+��f�1������dtp'� $��n��K~��$�e�u����rJ��<F�П��ғD=m�y|�*�������#;����|'����[{��)S�oN��n����Ɯ4d��^����'g���N�X�f��G�;��}On�(�����hJ��0"��� 3a3AA9�E�C���-3}�s�M��`0�m�u&J�U�T!����Q�����u>�Z�ƹ^(���d�*X���~k�:w뻹���P3��[����<D��Z����SE�=���g�W4��#��v�s��\@�)���}y�ݐ���n7k��^ʂ�h�㡼��<{�^pػ�9$�Y�V4�UEt<)�|�IM���R1ٹ��?Hhtxǁ�-a�}��P�o�|.��?\Yf��'�G�uw�������%����`��#����{��7ֲ�x�S�?��_ٔ:��pt�r��MH[{�e4�O7�)���
 /8�^�h�KG�e��^�XY�,���H���t�.�1�w����#�<�@�a��x3��{�qC»��Խ�:�)r1ɬ	�H��`,�	��#�I//2@وA<��M@����;�;5����2����Po��:� H��G#}M�]���M����3*+�Z�����Fȝc�am�J��I�h��|�� �u��OF�?��jg��t���`R�=e�d��1� ����9�X�/Q���?1��@�KeOnj�� tqZ�,O7扗�~��c5R1��}�,��/ ��Uû��!T7����T��	N��w������%\�%���5�	�p�_�Y�db	��JLe9a�\Y�5�$>���GVw�6���X o}�	LRdB���5��O\��5����#N��P�\��N�
&�/@l>��7k]AM���c����������=~5@��z�~��SVؖ�r2�/х�Ɂ�����x.re�sHf��]P: �Ϙy`މ��0���w:b0�/��	�b���&�c�K�,*��'�����
w����k�	T��\���{h��k����R$�r���֨�j6���ag��c<��IJCL��Jk)`�'͗N��t ��r�T���'����X?K������
��/��E�+\C�c��`�i�Sq0*�o�	+Q�:X����E ��=�����;�o������9��\(�xK��z��sP�Me_ϸFC�w�׍�/`�Z��3�M�����R�l���_�����:تk�h'[v ������}�U�/?k�X='�z9p�V\eX-���%Eؗ���QA���Rޑ��\�6���r�L����������������f���AvriZ-�v�R|���S�7�`�j`N*��Ȃ�V��Jl�J�4�T��נs0�џE}�7�ۣ\�4�O\��&�M?.��%�I�P��vЕz�>��b)<��˝J�Ň�e���G����	5���zR2i�0��KC2J7iz���Ĝ�Hѝ�Iu�e�/�!s���3��|�Vo�{h�1���w�^��D�}c��cn�q���\��&.�ȅx��?;Rg��'F��T���߮���,�<�4��;g��ַn�Y6���1��F�����_[݂Ľ��G�Ķ�Q3٦�#�>��̫���� �V����G�9D7L�l)��gb�K����/t��� a[���3nTg'�ǚ%2~����WX�`�FK#R�{&��r������/)v<,���|'j���]�t�]� ��3��^.�=�vkǀQC��ԓ��wox��k��6��d�{�����r$`���I��S�TU��c]I<O��.ԏ^�Dkq$)IC�Bh�sN@�@�'�%O5t���{�%�i(\W���[i��&��15{H��~�^��U�ys���4�_��t���s�w�j$�f��1�j�4�ϫ�n�����{��;ZO�%��&+�桃'q��I�/;�����U&Ax��}��[����H'K��A=�d��w
	Pk����:H�ni*���ZyCy h~^f���w�hK�vy�B���@!lCyP(�)'���)�X˙Îs��%9��/�� 4������HV$��|c�D7�U�W�1
@;s��3�`X�^����"���P�`ޯ)�i]�Vf4���ߡ��,AA�_b0��{'��}n����_	�1P��/c��$�e=q	E���e Y:��쨰?�$��3<�w,�[���M0�F��.Q"�˝'��"����4Ne����`7�0��3���N1�\��D���G�@M;O���;A)u�ڳ�	L������v6���*gGE׭0���YbL�65�B#Ӛ�k��S+; ��P����Ɖ��GU-/�M��!�.�o[�w�/�����DJ"rA��M.� �$h�b�_�J|�����8�͚F&X��`�E ����Tp��Q��1�le+��.f�-���_�K���/���խ��8�.&qC8�T�e2���QV��/���f.�k2ׂoˮ�̝�����k��lΞ]�����-�T߮��¥k��R'A�?��7��jLY_̖g��I��
T��`����e��iiP�U�vK6�'r^���{�]�b|��-~9qa���}%�©벏y*��EM���r�`+�0tZ�H�O�h!��a�����AE;!�]i�E
L��I-���0��d���xk�e���8�[~��䓕���
�W��z���`���U�~�xx��E��ߚ0V{�O$alLY��⬅�7.��5���Er�ӵ�-�Eq�0���:��� it�mޣ��aEF.LڸZ�W�q���S<z���)L��-�����i�� ���PQl����(��UM-��)V29��ou�(<|7�g0R��]���<�����!㰆�&���y����n��Y-d�!�4B���֡��t8��s�FAT#	P��(���uW����G��m����\���I�/x��n�x[Y`���e�����b�H'�.���|#�Y)c����:��2	~�Nl�(9�����[>�E��:��P���]��02�*JYU��{��t.K�0�1�1�|2m��G��C��L��9�x�Whz�!�K<h��Y|�<wh3���6����r?�r7���K���Z<�9I�~V����b�D%����	���?FVx�[(hL���<�m�u��Weҡ)Ŝ���N_y.R}xm�̖�{¬ZH�k�񗇞0E�ϻXX-�w�����G��l��G�{��Ý�;��`��^�������i
�/w b�[�J@+��q+�����zV�nS�Ʃ��
��1�A�q��S�5� C��k/�XՓ-��{ꭇ�o��q��\��s����q,��r�I��UZ�y�]2v��e!g�5���<����m�8�7d��X��qX;����}��|����ʍ ��L"	����^�O�����RY���zv�V������ ��N�65T��Ӆ �Qf�g�os΃��/ :����`�aC/䁗��M��������E�DD᝞s��!8GzS��!���IK��������Ǘ�hc$�צ9��a)\��c�a��Y��;.3n(�=u_ �oV��k�J�� ����|��nI�ذ��ܷ㙆�vn��;�c���� H![}O"\#}�u?B)��� �lok�.�L�`^N4�W�{���@�Hkq�2����xV�Dȹ RQ| &N�e�} $�I	 *0 �|$W�J�K+���@��ԝ��q�%�]PG���F�X�
�e�3L��48�,��"�yuB��>��^W1�]�/�5�
h���)�?��pi�o栽�ܤG��=��]�D@^c��ԥ;�>8��z��9�¥<	�ဲ�o�שv�i/�F.�+	]�O1 ���:/Kh�u�웳�h��ߌ�Ad�/7F*k��`Vӎd�t�=�N��3��k���;��ݱ0s�d~��YS��?z ��g���+�Kq8C���u�u�>�n�|l�c9V��Um���^�-q�F]Ӻ$�~���-���-5u9W��a�_��ً���Eݻ��:�L�_ ���A�as�!�OZ>�O�h&ֵ���d��V�^�D&�bh��+�0�#���^d����!C2�� �#'g>�N3qp7N:�S;�-�B�0�<TBFL�}v�p��]��I�ʷl�BE�0y���� h��Y ,�zJT��Oh�+����3<�4y�����i��=���T�ٮ��@]��H��rF/jih.���C�?ck�4��Q��X��fmt�Ks��lra��M�����J�X��B�(ZC��x�`�r^W��l~�$���CT�o�yz���.��m>	�IWS2 SzQ[i�[!M}]6���>U��6���(���XS�E�3dn��쯌
?�<@͡-��,��C�F��-�I��ۯGeɸ��Ҙ.���ȳ1�;-2BNP{TlAp�Is��0#`A㻢���p�-Ȉ�k����M�7�t4��P2	.Z��b	�䁯y�Y�A�Z	'[�]�?����F��\2	�н�t6��r.�BZOg� �/I|�W�~�o�c5�=����z�H(�c�K�� ���r��I\��m�U(r�d!�d�tOφő�O������:$�e�:���)Q�ȸ�&�,s��>19)�O��k�k����j*4�%�|>�l�E�8h�?�t��hzl<�{�UT��俠N%��[�1�=����ܯ�H�C���*���Ŝ���1�R�XDG%CM0���1��D�1��>�����p$A��J�=�CCS�H)��� ��{&]���%������lR"�=����8�BR��b�+��F'��U�ϴ�~��&T�%�q�����ع��*6�)��6��~Ӷ�Fo�K�;��'���X(Z�̠���V���g		�H3^�\E��p���t�{\������w�|5��,&[�'���t'"��╢gL��-J|��7`O������ٵ�;�@[9�nޭ���-�Ӻ�Q���B�t!�g[u�M2��m��bp��S�h!�TJ���~��L��G�A�cL��~���xB�K�D̃�x��$�����L�45W�Q�w�Ę���2�E��������P<����[�D�"�)�&}X���&����}�{��<����4��܅�;���rx��#0�Ȭ�-ʚ+���v�|]ZF�D����0��(Y���i�X1��<c��'$����?�^1oD��"�?�{P,DO�#�G,{5��H�3�no����U�0�a�xz|}���	cb��a�~^�$�� u�>�A��lh{}1Бm
�J)>��K���W�@��Z��p;Q��J�s������������I�9	9,%�n��,h���T�x��s?���/�Nt{6�|�Ɨ~�*H��W��ۤ����:9��Kp �K�4���k��E�)�^���?��t9Tڡ[7F�ԳXe�!�8�!�A�	�-�S�O6��3k�X�#2�W1f��8� �Di='�V+�a���gM��.��;)��N�6Z��Hd�E����/2{��:)�%<)��l-?C@/��ZW���Ws~M��kO�� ���ߴ��P��T,E�հh�E�Էٶ�DƠl������.j��~�O���C��s�x�.!��*�p��1L��c2.����Z��zt:�9��zuJ`��r����_�Is@kb�������؆�S��f�b6E��;Z�Z��qG�ᶩ����T�Sj��s%�/-IVi��cg��'�;~gx�f����'~�>^ч1�Ǻ��}
ؿ|�5����/��	�#�Z�Ԗ�A�v�C�⩐"iv8	��(P�$��uGD��I����v_a�HA���E|�X^���/2\{�4b#3�oći��Mf,c�:��-i,].C�_q��Dɤ.	ꥑA��Scɋ��0��>�2����x뵅���Ч���N~�U���[/T�v����6� 򍥤9� ���A3�[j2��cD���	I ��U6���P ��ً*c�L.���	5���� �ƻ��^J�IYI&J� �vc�՛��b��� /:A�Z���ײ��[�-��`�l�qh_Ym�6��#��)�89e�o��:Z��σ���Z�Y�=[*��9���L����j�W�R/�)�� %�;��)���B��̭?��I��yT7��]C�.RL9�3��)*�y�:�\��{� ��O�	���M�P�����[6G�4��P`&�z�q�ˤd*yn���6�|04>����Oze�z^�������2	��*�9֨��$$�}��z*�	$��ӊn��Z�c''p���?/��r@�<�TZ��Dk����n�`S��`M"�P��=1��G��Y6�j%T~�Dyߛ;�Z�v����/.:�eS��4�Gj�x��5��h��.�q��k��2����gG�tE�1�59<�+�-^�ɨ�N��,���u˽Y�n4xTڵy����V��B��ɹW���HK+"M�T���$�]����#p8p����� (KC�]ue�Jј~�\�M��kt��{����o�!3$x�"�~�ɚ�'Ζ�8_SQ�Bf�Y�����ex�rc����X\�¿�v�E���n�O`w���s�17���̼��(�+� _6�^gq�J��Ɓ'� 'J�sI�8�j�����M��'���,J�R�ߊ�^�x h^�|OƄ-�uT2,T��P�/3�ZCyOx��hz�1�?{�"/P��1��J����_k�H"�Ad��íjr8)?��[W�5�U�|u8��DT/_ɕQ�^�ÍA��Û�d�!��'���w�i�����w �C��)c�74p_��~�Zk��y��wl~�K
���op<2���vi$��a�s��1k}8|��� ��lG-db�䙍c�p�8M<�)�7p(�֓�Y4FN;0���z����F�6�7YZ;�����s�Ŋ�"g�#C���Qe��l6qfw�QE��Yd ��F�6�@�?k ɱ��@ж��J�u�^wGm��s�8�ny���nk�$����-�O�Q�FpVEl�-�G �f���hs�
��	��z��'&���MuX�@��2��X���}�y�����0�2�.ͲJL+h�{#O]-`�nr���3�U;SM�p����!�]���%2�h�vL2��  	��5om������P����~.����p��C*�J	(�/s1UR;��f�a�7�7/X
�Ŧ�[�r��/�T��bs�x?��-S�]rЋ�\������8\|_��$B>uA5=���{(��WU�tU.u���n���r >�?��f������]p�!@�Z����ќ���%Y�z��7P�t�n���CS(j�ytB����� qB��h��{( xl�\j���,�s��q�6L��]�Ԩ�#Y��7�h����`�m�������y�g��iY�Hy�T3�X�4��	�rMY�͕�����[�I*�a|~�Պ�N���]��IG�Jw���LN�J���.��?mx��1�X7�.J�8 �K�i���nϏAU�rĕ'k:��N��;'T��H��Ɲ虽��M� ���s�+9�x�L/5=�S�l1����X�M��	l~�(��r�X�1�'b��]��Ϝ�S�ؚ-9��	K}��_���π �_�n�$���"�/g�3�[�L^F0��YQ��TA�=x�#�v�5=�R��A�>�A��e?�tjn�Ècg�'ä,Xv�{�lb��������N���V���Y�ry�_!�Oz$���&�=��/��q*��'5:��|���d���g���<D��𛎖��y|�� �H F�P8zˌA�Q��8*{i�虗NP�wZӹ�'�E
O��#?%���$}8�2 �(��}�8�'�"lt�4��Wp�M���x�;��N�	�B8��j�u-0��6(B�u���R�nG|~֢6Ջ|�1���)�]�C�adl�1]+JM_i���$=�����zCV۰U�������a��"&a!����g,P%����a�'���0�0�/�7{z)�&���e�^%,��X�G
d7����t71���ݨ���ձ�L9��_��z44��GwDyz#��B�i��TS?\�F���r�ta0<�@��X(EB�VF�ۅAy�}+^��"5W���9�~M��\�̊_���
tϱ��l�Gt����^��3@�~+������v��MB�#�%}�5�n�0c)��w��:��mi�lS�Ln��:�T��;�97��V|Y`� ��|�����v��Z��?qc@����[�Kg����#�\���Pa�ZQ��������M��h1�ZE����#`����Z5vrB�Pn�뭂�J����?ܮm������N'r&�@�3>AG�ȶdC
]���{!���f��f!k��B8���DUA���b��T��bU�r��R<3/ԡ,��W��tI���l���1͉e�;��ž}4���;��"+q�E�!#��82ͪ�hD��8���D#�d��O;�D��gf�ׯO�
I��;-B���M����+>Q���0����0�~}�b��h�J��Cm���>���~CL0��@a��op]5b��P�&0@�9�9�ֵ��Źr�y�gr:�6.˓���\w��-�>�iͬ'���Z�*�DB��=�&s-3>	�c�l�{���9���!�|1�$���S	���2�c�;l�I���Clg���7�502�sx�oI��OuD����M��%�� K�6���K��⃱�8!7��ؙ�/����������8�P5�ƶ�g�������-������[�g���*�����m����3�/V/tm
y�,�)o���B�������+[�j�/��)ف7���\�������,Z��{�!^1ytm/"I���
��4���"	V8��dn��a�U��P��&="�uH�HG��o���dZ��|n��{�&,&���
 zDK_�J��W�mq�H�W��X�VG�WIB�Ъ�|wܠc~����N�5!m�Hנ~�\\�	l�J,��Y�&O���[��"�ʆ��@�!{�+:��$d�X�*�D����|k&�KA��b����9&��_ˁwk���OVYw��U�Rj&��X�l�4��}�C�H����.��.j�jw�%h��<k�-�T|6|�#L��@z�j��i�P��~�_T1��}f�g�ɖr��n�v=�?�S:Ȭ;6���-�aO�^j4�M��PI_S�O��1��V�#�>mڟ�����Ny�<;c�����|C�Lῥby�(њ�|W�\#ֹ��%��	�!8�F;�\���8�����g��� �JXғWPp�Π����Wx$�A�	`p}��7+&���0{�H�0�9.g7{��2��Gn�����Pv��:���]@;����d�y�\,��/S�����-�G����b6�&jk	�6��}��$5�_M����^l�.���%\Z�i�O��D%�>N�K �GZ�)�"��B�ּR-�u��^��fa�����%\ז�C"��k���t��AY�5����!�@!��3����������\� .A;��	�7�{cN�]��{	�,�Ϭ��í	��	v�.LC����51p�nnMᚋs�No��{��]��<��J��o�ӓ�[��%=C�9'$�hZ�=�U�*һ�m�␳�����B"Ŵ�י;�8߮�e�?Qs>V��8@�G5G���#��T7��1�����Z�q�pt.o�)����(.2\���FO��=��]M��)W��u��(�u�L�Xm�@�5!<��[f�0F4d���~�%�8+���B������|�H7�&.�43����[����*�#�v���܅���߶,�=��t��};�հ fu �,�#i�u��=�p��Y���C_�V�	烀���P���$@�:�SAB�R����(D/����&e�9|�Ggݢ�J���-�u�
OTL~�o!,�D�^q6���s�3)����[���v�E���ٌ�6S�ogq�������y*'#�W-�W	P˺�k�xV��MUӧ)P���biW��{Z�ey*<pA�q`�x�y�إ'!W�0pM,@.��~0F}1�n������A��ǯxI^~�R����4#;�����5v�'�B�uOh�O��I7��l���kD"�>�Ƴ�^��I$�w%2�}7���!��2|l�A'Hg����0�8o���:}+�� �{O�ϐ&�n����M��&��V��We��t.䅚;�Z�7�x�ؾ��Y)lK��8-T��: �O�����c[��8�\Ji�4x��͆�\h��9�!ձ!IO�[*�j��1�����sr·��=	'`���|ς��9��fr锒�겓�$�l^c��򏢞����T�9d����d�������k��i
G��R(hᔋ2չ���L����ß����jb������2���[��$JN8�Teh&�L(�kvȯ_�x
/G�"T����W��:�꼲�'5�*�'��ޑ�(t���� Ԯ��uwi��J�ФJ_���W4ֲ��~���/>��j$��i+����
�Sm�_��Cy�u��`V�	�jǏb#T��@Z�X_Y�]3�u&�å1�<�;���ȦWo��"8t�@��	4P-��B��Nz�u��h�,���ƈXh۷*�.}���u��)�[U b��}�/g��n��ؙ�0�waH@��~ȶ��Dh"��ݟw{I�l�f���T���dm%P�w�Y��С=��U���ֵ�K�@(=�.����%�&�,��6���;y�.�FV���j�jq�9G��"R(N��݅qm)����*Ư}���"�m� �Y.���_���7Q��q� Ec��,�N\�FRĶ~1����#�;9uP�Ϲn���_��yB-�p�͔�L�XCqaM�Y��]ϋ�KI^C���5���k��O�o�Bi�G���;�Y�{G�W�����D�!?/�s�~�	k,����+Za}��7���������D��Y��$�|S>�I����u?�X&ԥ1�N�w����};�I2��NN� n��P	��#�_K�	�8���x8��-�ڰ�)eJ;g�"��X���<�}
�T�d�~i�_J^k���Vy�ن	�d����!He�����uO�;��3G�a�=?�T���E-ib���N\�j��D]�G![i豵2���16���
 J�l8~Wp���D��C��L^oa�!u� kf�bUoy��s�l��D_ۣ���4�y�bpg=l8��Z��#䳢��\����7W�ހ���dE��f<ݞ}1���p�O�U�D����2t�/���j��5 @��;K����Y>��AY/�*\�+���=+ߝ�����-G�@|a�4�%M���rm�	|����ɫ���h̥��cu�!])�]�7�+�Z$x��|J�j�S��evh��D�ع��szj�^2���=������x	��f�L��]x�ʵ��*�j�����6T543�,��[����9�j(�Z�y�#%,A��D�6���s}�0�U�g�)>m�Xf�Zأ\�[(x:�ǐs�j���4�A�d�C]�^	�-�Ryp��71YQ��,2�>������>��")��ɾ\*�u��OGf��`�!G���>�ڱ2Uz��z�0��h��q���L�L-��.��gc���XR���:�����_�����Ne�����ٛ�%��S �]$e�C��޵�J��I,���̻�����O���� ]2�f�����t�߀OTڑ�L9��
�|:�'&��:�fr�k��6� V��iu0r��d�;o��RS�Y��E7q�-���BI{d=�w'�;ޚ�M��{������	*	;�0ı����
�,96P�jTh���4�&m��cP'��h�`��'	9H3����@	��G��J.�An�t~XG�j_����:O����/��Xw��ZH�H�}�q45	8��F�&`�� J�9&��I]}��q�Re7J����_D���
��r��jE0�h���=�j�޾g����8���=�D���V���&�z���^|te����JH- �����^xخ@��D���A�h�#WT��'H(��x��k�c'�y0�K���jN-c�{28y�M�ߑ�v(Fs(��zF���m5.j@P�a
@�]Сp�G�	hY�)�X�dh�-��l{���۪�����O���O����ҟ�Y�r������qX�}B%��2��#�8C*D3E�"Dd��f�ng����%��"�O�2����JW���WxA`"�i_���ݰ��{�����;�K(��>�����_�T����&l&'ā�W�5�7���rY��烦_��K��^}7<C"Z����ռz�~4�\af#�$���!��i[·o�/��.D@Ku9��]A�\������݄))O� �N$��z\
A\�W42h ���4�!U�f3�z!��U�u������{S�C���ň0��������5p
=��i��$@�� �3�M�Q�cɞ���Ј\G����"�r
�� ����.ϻ{u�l�*r�ae�Q	��wG�ԃ��V]�g��m�Z�w�zBc_q��V�'A�GO׶�,ŷ߼�T��
?��m u�G��$��S��3����&PnV (�@����@m��1�;1�{Y>4hT!�Gk���?�~�3��䨩�[�U�̇o��cy\ �������G\ꟓß2S�R#�p�n�/��h��C�XC���ّ��-����z�е�&'�{�TH���'�����{���B,;VG�H��������:_�-m��Ur,|&�N3(w�M=��Q2�`��J�ج�Bw؝���7�Q5��^V3>�<�XSRx�!����#����*^0�y�
6_�/k�m����V��o�lh��.�kg�"� �y-�w&���"̳
�=�i��	*��v�� ��[cX�9-�` 0ɻ�����Yj��H�Vc�F�B,�;[O2BIM=�k�g�p��H�V�+;��'0���γOJ^T�=<�=y�ޟV]8Z�P��5��G�i~��ϔ� %ua��:��.�y�t&�k�\Y`G��8opA�x�J�� r�*�t�<i�|e)�ϖS���*pu>y�+��i;�}�Z���<R:�y�>��s�ޙA��Db�s��O�`,�,�_X���{FAk�����vy��2�o�|i%�2���M����Ũ�O������e��aZ��uN�@M��lh��{�Պ_�/Y!DI*۶�̒\��u��l.AL��R���°�ߞ}��^��io�Q������QC�Be4V�E�e��C�4��3�!Q��e���V��Ѥ�B�y]��#8.���^�.=��--��b�CЍ{�9V@�fz�:>S���0�޹h����NR�{�;��<2u��_�V
%jԣ:��)ǝ�sIXg���'���}�DI&�l4��Z���u��$&�%��72z�0�c\R�O�0m���kIExB�Q@��9䒑���^I�0�9
e��;�o���c�n9YE��H��P�5���<ۭn���;�����ft����W�j�^�:�2)u����0�A��9A�(DV��v+DĤ2�|��vhdE@..Z�Y's��JU$!o}̈$5� ��w|���Rqę��+����4���w�ai��>w&G.��T��c����W��z_�S��*@�2��5]ȕS�'Mn}�zR�~0��Ho�W��HE�w�`���yn2B����:]�]O��h���������8�f���"��(�mP:�ŅQ�F�N�Ѽ&�!�H�"P�p(��ܥ�����g|�\"2W�@��j0$�Ź��G�q��t�_,��*٤?�`7�J�ea
��k�3E�o�: $gF ۄec�LN�Q�F���o��~�h�]Z�9Ӻ�k �P7�}\���f��%�H��lH5��/::��!&@{I08LX �51�㟘9w���@�BEk���6F���*U�m�@���b��=�{��kŏ��Sb�2��w�Oj���������Ί�[6N �^�Q�=��(�z!�M �=yv۲�����YOt�ŸTT���:>�)���,��'p�o�Q.<�;3o�2�����a6~�]��D���Z�wU'�mZ3���ᩡN	�@K�����`� i�N�Z��v�5 T�8��L̟	�$����:�c�����Ga.��� �Y]����1���p�='AQ�a�0����_��B��W�����T�]��8�bN��YJ�b�+��P]4r�F~��<Z6�����C��s�`��f�z����H��'ղ���3D#���he�(eЏY��l���exY1�������ٶ�g[�ܝnd�5��nS>0;y��`�hAd<��=f���4�[ �J�\�߅�E���hq{M���:��+OP0�ʨ���L�S��L%u_u�  g?ȴ=H�h�I�c���叢߻�Ŕ��$�@�3K��k^/�S�'����NL��
N�{Ք]lz�:��є�~euN���o_aF�6wK�m��*A+���쬔��?�X�I�h�qğ�}�s}�ZE+A$g3b�6���T�
��cE�3��5�P�� �SX�n��Շ�� �I�E����-igH�ϼYE(MR]s*�cV�:���ёPW���S����R�ؒ�1:&���d�+Ry�
�w@_�n�;@��T4�B�!��$�A��v����&R U. 5	���ݖ��Mdlo�����<{H���.��9-����o���l��5?�5]��C����^v8��ږ�}v���ʖh��v�$�C�ʐW0��'M������- "���365���gͶ�r{^Zm��[����X&��M08-,}��W��R�M>]��dE�*V�B"��H�^)eR7�9Ε�1c	����,�� ��d�����WHq�HLDC�Z�5���i� ��rvv���<J�<�T����tA�E�]7��3��)G��;�3';�U�uTU��IϪh���P�o+|���L���i�T�z �u�U������U���Ol���~�Z�l|���W:���8��'E@��./B��������[�a� �Gm�9���<!�ݡ(�p�u{Фn�10l��?{g\�����e1���ᗩ�(����Y�H�&n�7f����J�(�|v�"5qy<���qk�xR*�o����K����1�4���B�����u�6�/7.�5%��0�]�'�d^��8�9F�����*���<�P�HHd R�� �Fj�
z"��,�qr������4��Ě(t��j�4�ѺC��;&�]�P��ʩU7��w�x2A=���ܾ���ͽ�3?��17�ǫ�)�QI��^Z�H���#�+Q��a��n`�w)Xǋ�e���e�����E�g5 	�a3��5G�k?
(�3��9T�2��ܭ�[��[�SBb	d��3ɞ�� �yЋ�kQG@Ӻo����-����KsQ��|-�ʌ	,ޅ*���2d�8��R�����}�(5����%�]�v���;$�EP��.��k�,dC���$T8�&2���?�����#r|'��#B�_� �����I��8�K�C�z�M����<Ž�����ߒ�B`��i����5�K�N��,iZ��K��+��N��Y ��IaI��\�ٺt���%��-� ,)��\a�ѹ���0����.#��>#B�r��3�ߠ�ۋ2��O���+cd3�sf˜_2�B�#}�TCbCSeɻ�X�<���i�ɱ95��#Cg����H��x���6n�9�X�#�P,����QO�����a�R�q��[a�~hB�)�����[#�`>u4�xq���,�^�r�����i):i����{J�b�XlW��A���_��f9M�;.V�4������G���*R���m�=~�u�Ffe�������_�&쩼1\�%��3�y�$��%��oC��!�lƴ�lK����L���G�
��T�ϱמ�½�I+�՞�4��_�/Mj[��Q��U@���l�A��E���E^� ���
��)Mn�Z��(
<MG�WuPڈ�9����;���1�_D{o��s����5�LO�����	�$�����w2��5��d<}��[���/{��7��p�uz�D��>Dby��@��TI-����~FeDU?)�
	�*Үqjg\�W�H������*�������\	L�Mi���Fs��Pi�F^����b�C6)����-��u�r���3	K3v��_�����3������ZNB��~��z /�d䙉����qJ�m>��T��iv�	��C�Uܧ��r|�\UXؽP/��-����Y-� A��x=�����+�H���$��p:�Sȹ}OM�q�"�Am�ʂt�u�w������R�yǲT�-��#M��} Y�s#��ϫ�P����{a-�m�O���� Q����sa=R#6T8�G���>,�#�eY���E���΅{u�U���F�ټQ�e,��ܱ1�ݹf�.��(-�u��:#�[��_�lW.qT^sO��V�h�:m�z�N�;�4+��ҧ�e�7�ػi#B��q5b'�{f��!(0*	ţe���
}�u�DQ�rs��^i��Z�&���pr��j�rz��=�<�1��I���+6>Ɨ���s�;��,�KTS|F�R�PMI�+�q�~��v;gf����^�>�8M���C�U�2ޣo),��,>�7���~"Hi��\��Վ��?H�����G �p�\��6
�\JǊG�Y�����c��^r���,IFh*>���lg8=��w���� ��o���!'p�7�e��bq5WIL��a�V܋.~f<��>��VP�Ptv�E����u���bYg38�72\X��
��./KP�P��Z��YG�A�h�h�Ȏ5�����؜~��U�R��VRH���:-�:�0m�lRy߮��z�cÑ�Fr��, ٌ<ℾn�ٳ�-�}��
*)�̾�.�o��a�Z���%��s蔱���G_��ʥl۰~^P���Q�mе��ν,�ۜ��]�k���A1Z�A��,�[�C��?��]G9j�75�"L��n ��|Bƈ���]���D�6��	�:%��q�8nZ?bj��a7�{��{�9����ׁW����j��mq�;T�����O-1���~�l�����4i�aAgE_��ȨN��Ȃ���h�gJ 8g�_��XȬ�>*�E�;4�Hޘ� �8w��0��	
�����T,	n�B;��2�_�#h�D�X�g���#�bDd|���
x�EZi�ޑh����f@m&n��l
5���cL���r*���V���$�}*S��u�ɸ��6I\02e*&� ���a��4<�A��<K��w�꓾�!�,��c�dW��@u]�8$��=�E6E�HN�w^��{�`۵����?�N�HP7��Z*�Y~�̮�k���7��!���l�Pxe�����e,�l�=�� �K;�н�-Z|K���X��p4�wO�+#�E�u)���t!�>��[9+�,�`ì���<���{ƪ�B��9w��)]��b��g����^���B�u�&�b����=Ǩ��$x��Ț�F2ە��/o�@j�_갮P�t1ûm�2���_4Xƞ�c`��ˣ�	�W�~=��Z�+$^��,i�]� �ܕ'�o���;1�7��:#*���h|�F�&�w�g}��&pB"�0������n6VQ��5[�h	_B��TCJ�~K5Bd5i�<o�Z������ǡZl^1����Q�/��Ɵ�2:�$`Jt�.�+C�����YT�?ܙ�E��}�ɏ:�����[YK6j�/�	��@%����W��H�<]�6_��~o�?6/���F�����\1���P>0�e��H(�<���L��74l�l%�X��J�ُO��!�L��U��T!�M(`�ry��#��j���ҴT��T�Ct<k�o����?O��P�v�0�oҤ���HǤ�������{!�'��ʷw�d�r�����ۉ��!�����~�{���i>�B\)�v�b�[��{d�J�R���%�M�}"�����k.��p��9�K�F��Ѹ�_x{]�Jn�L^��h\Y�oM�����m?��9A�E:꾜��H��^�������;�q�T���qS��y���ع�27o��_DL�+��;���ȍ
�c6!��0�E��`�
��Q�HGۇ:N[�x'R�)���F/3M~��Ï4c�j#TkWEȧqߝ��ګB1E��D>�~�:�����Z!8�A�4`a'Ǭ�&:��o��9,k�d�1�n�"ND��8�t�r+8CIҘ/�9�g�!��<\2��]����ɕ}���(:�h���Hu��*p����<?����=�s�\�e�0D������P�&�5;p�,�MD78�~Bc؄#7��^�+[���>�]�N�pɊGI6�:�Ѣ�@�����i��qY*�}Wg�@�� u	. c�^���E����V�a0~���H���T��ᥑ�w��-aKo�q�~D�t"��g�m=�������Ӏ�ٓn7SO�������7�
�y%��D�WO��̀A���\���>��ʊ �8���np:��Gw�@�	I�&��e��"�c� !K�#:b�\-L Jv>ʕy���z@W���U������	����;0�u�6��e?ps���L��LW�P}P���/�.l�D}�.�g�M���.1�o��(�8\A��I���Zx��?g
vx���i�i'+�)u�=�h|����q3�����~��U��~�GD�0ח���Qv���J�7�x������5�,|�UƔ�X;K�`iK������k��Bmx��u?��`�L���@ a�{9�	"�N�E"W9���*��^�v���g�PT��A��Dԏ�10rC
~!w��%#� �C�߶��/s��E��l1-��;Q5�MZ�@�4x�a�9w>�8c ǻ�8eIp�T/w��Q��᳅��{�9}����\"��@���J�dh�U��	(�AH���dg[o�Z\�M������0���-I9�p�`70�G���	�<p��N�V��K�C���4�㕐����Ȕ��Wά���̺\6GR��)�ˇ("d�d�l�I���͍��߂l�G���И#}R��i���2�����!���rR2>/R���D��ޣ]9S�2� �z&i���O��6-��f�2i�Y�_�u���Lc
u
A��c?������3	��Y�����2/�<K��Q��dG��Ta�"xEH2�|]�(}x�����z�/�UJh���j����?�����̌x
���4KP qh�C�_�p�'ƹr���P�zz˚�|��G��,����6��_{�t�����yŇXeKf*�������X��g���D-��I@��F�E�$�>�7�[�����^����ΡK���������[�2z�Mu���lb몇*��U`�Q>��mS�șm]��EA��UQG�0�c�������5��K��	r��3�ǻ\�Zr{�.{�Is���?TH�`�Ѷ����\����i���!P맫�ʪ��c8�k��M�4O+�P��^���H(R_⃟��2����{惎ȃ.��R�&$��C���w@��V�Y�'gM~wp�x�R�1�3�׉�YP!V-�&tN���a��Mc���"������aX�)�������1I�)��ƛ�S��~s�9睇��9�zSE��J8��ly>�}P�a�G��t�Y�r��vJ:�Ʉ�x�����)t\�h�ޒ�;����&������N�$^�P,ICkZ�M�` ������lɯ���h�y'㸃"���D�6���7:�Q�.G��ڷ˦M2أg��
�`��>X�q�D�д�˄���IPƞ��* Y/<}[��./(��48�2�����|��1R����1�I�&X�{��Fv��P �t�0�Mzq���������H:�v:P7b��A`9޵�Z��Gi�Mf��Pn�2���ڈew�;�÷���/�O���P�����
?��c�o�b	{IH����o�sO��1�)\�#��b���[j2�o!�����v�L~�O"�k½dj�1�`�-'�E��V =b)� �m�[���.��\�#��L��' �0�! �5d�Y-3�Ίa��6������Sd�S�k���Hz��a���[�_��u�O��ٜ�~�_���Z�����kSSJ�r���|��/Q�@Ķ�,�ɵI�Vs�שޑY���:�Բ����!��+e�?|�����=���Y*I�4�O��&~�y3�٥�\w�{�N��L���b�M����=O'!��m�S�����7s#8CQem��,|S���Ɉ��6��#��{�����w�8o�&�/���D�H�j��.���Ɛ���.�5G1� �#| ��æ���Ƿ��ЎՊ�[���ce簆+��i{�+e$�b���̡�4}�KOg��bᷴt8��I�tB�ˀ�}a3dy\M	^8[�5~)�@2�h��X��QvXD�jD��O���t�eR�;�g,�QW��q�gSD5�I�[p~������7]����f��Gխ6�J�2 �����GN�:�Q4�YoR�9�3�%bu�t+������4��ڸ�t8�������r%Y�o>��c�!��D��k2C�	�䲕�Vt�Ȝ:!��佧g��`V>�	��b�}���o�Ɂ�s�"�k�r����-h��J#�9�ox�R�RυŤ���Aj������s���Ø����;B�����:;�������k-c]צ�c-*�A]:���ԟ,g��K*�!g�i84�,���Q��Dq���W`SO���!�l���Z0�d��aޥ�����+�K%*�	�$�
�X�	�j���n�����������?�3�,�nY�=�9��Eڍ�xGهnKj]`o�4G�ӹSG6�M�И�>	�\k
�,����U	���� Y��~К����^�-��ᤣ�C�u���C�J��j)A����T�7u�*�f`��a��N3`Y���{�3<�"�Q��G�s*[7T ���ޤ-H���}��;��o�g��������1s	J��dmK�n��s'{;2�d�O�{�:ed���2�%�%�͍ß�r/FěZ+�J�����L{�#�t���o�韧��\1��F"�m��GH��rz"�+��nJ&]�g�?�l�8�_s��I:'*��.oFtq�����o2�%�iă��I�M�J�	��wq�������1$Liz~�8�4��s��+�Yt����/b�H�B��θ�p��.?�i +Ǘ ���S{��"	)��;�NQ©p����yA���tE��r�
�C�tőF�+K���a���{V�Ҕ���j9
�B�E"U�t��G�
㳤��GzB4&�s})��dTӽ�)~�vO�r{���,����uk��a*�fϣ;jͲ�1\�{y���䩚�߯Sq�v��8S��%9R��Ĝ��N$�Ȯ(�eF�>7�D�AެQt��gqL���3LR@�g�^HȤ�Nj�^��+�6��
����x��b���`��f}�BN��=Zn�v�����nXe�srx�EZ���Z�.����_����?�=��A�[D��ȩ�W�0��6�)q.�u�W��1���ƅs��Jk��x�ԑ5�DsXaU�Hx)w1ʶ*�R�.St��5`���]�ug���̕T�"���ȹ:�0��O���^*.�}��Ot���T�?hJ�[Wt>(�#u�Y"�gT��P,y_Qܱb��Z\��tJ..��;�b�"h�!-�WJ]���o��~&]{8/ҝrg�����o�R��s�����i!ɼ�������Ȓ����ż���\-��Z��V#�wpq3�����9҅�r+�ѩYQR��P�wo��є��4��N��.s��g�8OOs�в�ͭuq�"k�~|h������-���Ϗ�
M@�^V�U_;"|��]Qɰ4���_rͳ�y*����6�G�(�?���9�2�311~�EjL��3;C����������
�>�c������u���c`Zr���`	!�
�*Y�f���C�ly�p ��t�j�`G3�)�V+��%3�-�}H���S<�X� -�>�:͏O�}�+~{5X�b(L��9�u"���߉KB+U���Vud���/���o�L[Cǿӵ����_����"1HI������Wj�BI���S��9���kט�T��Ֆ� [W�A���4� u;�jB��IPռ�a�� /:����?P�P�k�p�;���� Ki/tx�|?u�ԖZbL���x:�S2�E���cA����6�<�����O�JS\o�m��Q~C}�K����z3o�yv��ye2���>f�f1�_��F^By���1���{K�V&���jj>:��G����E@�]<)6�����&�����Y +2���#`�Wu�d�������p��玜�)��B_F�X/��Qp9��#�L���l�k Bv��$�U�(�]�$�V���/����ࢱj%��ӝ�n�2��1��d����Ϩ���a�L{��v�:X�O����]���T-�/�H��)�:7�/V�� �ȴp�Ƈ�O��U?^�"�?9 �����C����ʿ���^����jԞ�Ƨ�R��l	���:Qn���ׂd���"�8;���n��vZ/	�%p��g�E4��-_����"�R�8� G�rl��X6�H�ZМ���B�aa�бT�K2�lK)�z���Q�5|�;:h�:��Y�Y
���� ������!D\f�z&�TQlS!�_	�	���z:����=�˨�MC	-bv��w��2�"Y	
�	��Er�ə���z�Y`����8��v��Kɝު'H��1���ħ�����I�Ҩ�,Z&Wў��[{��F<#��Β�S�J$�F��� �`�ȭ�2S_ SeO���*Z���9��'bM�Kʚ��U|�����d�����N��Ʈ9o�Lp���窋��:ڵ^3�:�B[���aYD���*:8{P���P �ޡ��K�W" q�����oس(ѝѫ�6Mn
�O5l�y;&���Wc���L���@���������ƍ�0��Y���b��Q�-3�Z$F���ц�<��8�Q�l�-��a��b-�fUN��a�0W߳qd�u����z�)0I}aɵ�Na���<ؚ�5���~����!��k��-t���k��A�5U���R�G�l$��6��N��7Y{v��R��"A���f���\�)�'h���k��D�����[��[	���ˆ��/��,�X��{��0e�K+��-�� ��6���e��ՄϽZ�U��$�����'U��S��:�=���U�:��W^n��S��>ܢ�d�;ؓ���.^c�G@�)8�!�&�wL-V=�D�=��aD�7'ʴ������� Q�!�K�82C�n/Һ|����!G!3��.f��<Y�~�⋟?( p��~�u^b�g�j$w�?u��t�k��㑅������y���krռ�!����P�������±� �� ���f����뗕������{��WE�x�&�����v�5�]�;�*`���z��:��T����etY}AM���1�Y�4ܵ��\,Ղp���+�]�(?f��U�Y^'����c��U�� �P|э �AX݂�א0�־
��@��i���#����� �gIPr냕x�~SoҼU��INp#v�K݇Ӻ�ះ�u;��������|��.�zөG�¦�.�����ŚW)�7�&��>v |[ƨ��U�]HC[���7l���������C8���I#Z�6�hh�%�N������Ɇ���`�d���V��=�@2B�j�/�;ˍKڍ����ʓ5�KGD~z���%H-�gA�5�r:�;h��a�n/1��аwtAn��b�ʶ�;�YӰ�H9!����4��/�/[E�`Zk���g��$-f��%���b8hVj".y�;��!��G��'��EK��DM�0t�J�h�M�	�� l oD��Ys'��z���dP)U��_�?Zn}��).AF���>9��cM��}��a�j�����i��8�x��QW1���UD�H�Q��b�L0�bT��[�7������,�MBw2����^������܏�%.���X�)�,G"$40�3�P!s�D��6��<�M�����@u�z���y���8v�/X�_��P�lI{�4+c�� 9F��T�ԑ!�xS�l=�8�#�=�ޭ~v���&XB���\�u�W�rV/`�={PF���% YW�~���#�G)�Fy�'�j��\v8e��I��J�����A�4�ݧ��ɆJ��ˤ<?]c��Xt������p.l��h(���sh���P�K�c�-j�߅�\���C��1�4� g]V 3�:U:H,�wb;>c�ɠ�F�),ѥ�_0�Hf�c�L�q�7�Ϲѥ�_@�b���	(�i��7�%`1�q Љzc�Ѡ���	��x��%#JedQ�YMNE왅����Y�;\���~�T �@w�S���B;5���sQ��K�<�A�C
�$��Aò|r��q�Bh-�M3xH x�5�l��C���C�ԝ�r��v��7:UPAy�I��{��[�?̘$�C#ܢvTn��� $nM�T%�'*W� ��	%����H����(Q5_�*9gˢ{�i�U�-�9����"�N��ħB���X���A��y��8�2 o��V+
���Sl�vֵ��[a�;>����p�n3�
~(���T�܊@d����8k�F���&o!_A���)q	s�� f\ryޛ��j\�*�n]��/��|��-G�� 9 `�R9}u )����$f��O�f��� ]�޹�~�����١0�3�.��k���ak�#�I8@�#,�T0�M�i\��TYW�{w'Ђ�pV]�LJ'C�EK;�/�T_�i����/������::tYy�"�
���T�}��8n�i�_D7k,g��*�����O������k�EqY�3�j�L�>��u������^saK�@�"]՟�x�
/#hM �G�N��!,Y(kKb��F'� �1]o�M��']et*X~�1}���[h���3�����[��ɖ	k�F�x5�#��Ӧ6�(�V� R�;$)$�ӻ ��B�5%���;�g^ܯ�T ��D�f^~S��$E��o�,|��"=����&��wq<�������� '+X���9�:��-|����0�Vʆ��H�ƫ�$8�X�/h�8V��<��b�=�j�}��ULY�-s��Ws(�B�����Z�J��*|��Y��z�g>�:��bKL\����ai�m�tD
2AtڙWyb��EiZ�`}�}E~���T
'�_0���J3�fȁ���6�y���/�{���U��N��X�̞���2�cڱ��o��f�Ą�m�547���R���:�[J�L2�_���-��`��ލ�۷�a!!�1f�o���w�2��=���.�����P�H�N�s#�\]joc$'42/>˔tN�q��%ǈ�D������r�X��䶫���{��ON�����Oq�e9���=5���z�f����e���nu���<J���\O�Z���:Q��tw&'�L���c�3���(�����p�����čirhQ��Knv��ó��\���+-mBo��6#
�c�,��3�b3�N���D�AzUb��_����{!�����\H���klgx��Y�r�P�%��{i����'#��&
!���7��0E��1����7[f��X�\��#靧
��W�oQ�����,��0����B*p��d�S��-��pyc��{����g6zM��E���
P�Fds=q��P��5Ɯ8f��;����e+�4�vFC��c�/m8�g�q��0o=\�`*�J|gQձ��3J{It�_ H��b���ׅ�b��f�g��K
<�*n����3�) ����`���4��Xv�^�#)1q��+0���X���Md~�'x˒�Q%܌�g��9���n0v�ː?>^���Kwb�h�Ͷ�a����ͷ�f�}�`��kS']�⃇�I��s-��E��=�B�97�j=/0��.|��7��Riη�������٦��IYp�A���[ۛ�BһU�1��MQ��-H��_����9��O�D��,I�Rq�]����I,�a$ONw �����X/�QAvvh�0���ǀ\w���Y��7�H��O7;��D�ȯT���q��jgpt��������"���|B�	�E����0[+6D����g�ҍ���|� �&C߷�{	������{XV�Ԅw��
�����K5���n�����u�<�dmV|�0�鳉 �e�0�j'������27bM|�j�5�T�6Y�]5vH���
��%m�tŤ���j�G���ml�����Qߕ�XR~M�K W�hfS����U!0V�;i���42��->�d���!�&�,�s-B<�_��!���������'C��6��gȆV��O�AQ0�X�I�t� �0&�y[H;!�	�vъ�Y��y�+.��p�e��Q<V��Oo"�On~|�)%��{-0غ���7�����aגa����뱬�D=QJ���B����-�s.߱���I��y��hv���~[8�;S v���`��ց285��ͯ>�K;H<&y�5'�5�E ��Dӛ`4lA���r���L��N�=��l���P��N�����kV�_{
��{H���).���ʂ�#��I���$��lF��JD�-`(����D)�7�WR�ZR�c�jA�xt��
#Y�_*��oL�yDy�άy�N���r��=U����a�ۭ�
G����M�
��P�xa&���'�%�ix�zCS�͛g`Eb�W���5�<N�~�s��X���0��|\�bU� ��0yI�
���d!���Ar����t��B�'���'IE5����ǆL6�d����G#��K�3.���5ҬB���-���,���{��q��G� ���t�M��v���&�P!���W�{�~�59���0�@;~+�kz���ig^^zs&;�з�;�IKL�>���!��	��N�gh�t���5
�-\�4O������8�>N-��)������J�ש$5U��e��_瓟F�L�cCH�Iύ���cEf���Ժ6V�~���v����W2�9��]��{B�q��7���ղ������NiQ�h��ch���V��O�cݤĽ"^	����!6�t{Ǌ�1��C�J��ȍ���;2��T��t9��e��sѐP�Xfe�������ɬ�P�����+l�,��?��+��|�H�(��3��X?���ĭԼ/n6u�A���W:�ư�|6R�����ޘc�%�����F��/�>a!!�R�M���VʯR����M!E��vJ4q=�@�g�44*wG��XY�a]Q��>�)�׶��-jX��&>:�0b���Zd`D�t�!�i�O�q�lƾ\�X:ay�#e�ԗ[iǏY��Xݤh��lI<�}m�iJW$�7�����FMj��2�����yĉ���z��j?��J�un.�P�; &�i�0�ҦX{�[�C�0PJԃp�_VO���]�ql�at��-M'��3�ZiAo&��[�B8�����\�	>�mF���]��|�̙�m:�s�x�GQ������4K��  ����Tfz%n��+ArsI������;�L�iݪA������:,�٣�Q�P�+�X@��r��d���̪,��I.���zMی�aY
�,G�eT�a����w����+��淩d��|���lK_��Ȣ�{�R�����TUE��q��q�1�����2��������u���䀦e�	�%t��(���J��*=� C���Z,"�kS�k��}��ؓX�����52I��
�Hz�(�3���K�����ovJs�Fa�æ����fkC@j�vUd������d��[H� �b�i�do�Mi���;*~�5�a?��)����'��I</�����n됵�U����O�"���+�amd�~�"C3ܶ#�����j��*^�̙c�0�Z��̠�A�sC��I���`����1�e�͏2�S�Ic��M1c22��qK0��`@^��q�\MA��[���&L����'�5�rm�r�'��ύ�>�2�V��I �p�2I��?��f���,*��7]A�>����8��U�V��`n�d�W�h��E���@�9#s�bxC͂9�{&�O>��EV�i��H�:ѠRZ��;NRW��Ԉ\��-e���rV�1��Gjz,��iH�	N�N5�Ð��0�Y�����y@&6z������#�6�#�F�j���z�D��\�����R�T'n�Z�8"�\���,�@�7�`x����Ž���ͳ�)l2[���T12zr��A @���@�߿��������q�������/�6��
M�L��	�0�v`�C����O�]�1��@Ɍ��>�k����>e�F���/̊�rbdHB��R9~;�qn(�s�C����D���\�Lo��[�V�Hj����u,ߛ'�:���ˊ���R<	#�!��t���U��G񜟣膨���EVփ��"G��쓰�����"(�6ˠ�n�n�O��(���Y<z�t˜�"wL�VNL�+��t;����x����li�����r �)>��9j�P���#;&���sC�c�:��0��񄀸A}�A�\�E��
Y�j0��s˹v;��2�:��E�}��Nf��e�4d�����La��YB�������0m��H�n�X��^��P��
W}]���½ר5���מφ���h ��k�y������3T|Y ��POĆ�����cT/)g� �xS���fy���$8�n����ƽޱ"T@�;aa������A\�]������ޮ�'�J�
sc�@I�_~q���	�e \_aR�ֱ�a(�������w��C������%�U��7C::��$�r�s��MXx�n6�����b;�Z��;��m)����oKD�MgG��Q`v�9*�Q��p9&)/,�s���kO�K��k!@�I���L
�y�m��'z�Ƨ��^�>mg�^pԵ��=����{��7*N{X�\J�� ���?���� �=`�'o�
Bg.�2���ɖ_��T_�ӱ���A7�~7�)J�>&�7�Yy���C�?#�ׄ�=��{C� ��t��3
W@%`�����c1���;0��R۱��o �J3�@
�r/��4f�~vߖ2#�\�5�u��q�M�[	�ƣ0_{���k�Z���0ɥ	�
� �x�RA ��E��c��7�jw�z	}&�$���_���I
����Svv����w�=�Q�c�#M���\f��i����oJ��j�w��0+�^{$��/@ǰ����k��vi4�k�9�Ll�X��=�g���7tG([|ـ���T��9���3��B���A���聀̓��c���i7�����8�&�9���9]�D��;L����R�*��@^;�D�s� }o�8��\������������ҧN^#�����Y���<?['�k)t"�>fY�
�x�Ѫ�@\�K���i�g��a�C;�ʤ�HK�%� �}�����(:�v�تB�9�YT/@���?q�N5�ma����R��2ˑ� !���z�u����M'�6��K����_TL��U�CM9���tj��H�Ut��	���5'wu�׵X[�2TF��T�:c&p�Q8��wW�.;;���3\?=y.T�R KH�ҝ�62S���C��Lᳮ+6#mmq�9�b�3w�W�Mr�����?�z��T�!�<�H3�)�T�+��m�M������<����?U���GH����Mdu<���H�_���w�C��0���h.��n�v��LK����̅21&K�u<`�ͨ\�^�P+%O��d��Ĩ!���6$�4��Bڧ����X�%$�w���zD��סxɺ\44uy��W{|�Ҋ��d����m6Jb�;qp/�ִZ:��Q��1'D��`��~|9��������!k�CJ��������T�!k���unfR��ڨ��!�q2<�|g$`�L �0�xL�Y_�& S�6r�;�@�8��@Dd`̩��i�
���;���-j�5�A�L!f�C���%1���;��)?ev\5�#���K�V�1�d���=y~ɥ�L���j`�0c���:���X��\,�RY<*>�X�(@��zg
�l���&9�U���@$x��pJ��@�Ȭ�G��C��eT���p(2��H��W���d�:�QHa'Yv1��p�l��y��x��ѩ5����N��žX�*��.
��(�0�{)�s�\r�3�ZHl/'� �>A��׼�Z=`����S G�&��.���>�?��\��~5���MBb�I���ؕy;��|�-�L���y�\����nc���}K�Q+!��`��Dy�D��	Zw�3��b�#	
�]��Z�o0����_��:�Ὧ�3}V|Ԡ�|e1�[���h;�̣�ۣo��ʇ��Ng��_}��5�[f��(̃b͐�B|l�0p����{� ]e���wDwEY���o[���������z�	� Z:��"}� �6���k�ӯ�Y�
�$����Θ��0���F[@��l���vP�r�h��σk>8�XrA_To'ȩ�"�	�h�%��6W�˃�v��!me�,��SgM>��N�/���[�.�Ouȴ����Bc1� pΔM���h���k�������:K�n�d¦vl{J��$�~@���Cn
!��?f[�8�vP�z��7�&;s}���i[�>e"�m�>�h߮���>13����r8Y��"A�>3.`O��z�nvt�g�=�}mW��I���:o��2H�w{$������\O ��g{bwQ�*��6��F���t��Ә�x���#�3����<r[��x[�����%���[�	ʺ�L�έ�y��b'-��)��d�v��C���ǎ[����21C���L�q$�
$/�`���\���Cm�8��F�iܦphۂ�%�Lt}k@9�E켫�O�ɨ̌�yǃ�@�B�J�$�^t�I��^��R�鑁��
�� *��e,N�D;�w��4V��.���r������B)��]uDO��z5G�9�>-����O>�}���K=�?1����Y͹J�tN�!: �4� &���@��+�˧��q�1��x4�&`�&���
�Q9��G��p-4*��?�
W��ʨ֜%��1~�Q�+{�>�?h�R 0(�\l��7��O�������Ӡ^=����l:5A��*����7y�Y�>����Uw�Q�~�����U�޲����h7=�@K��~��{@�MНI��Y+i���ȳ��<,o��"�T-�NM�0x�=]�ȓ�-ku=����"�~'0�C�<aѩ��|�A�����=9h���*u}�s�"9Ek~1pmb;j�x�k���`Z.6Z�������MR�K���iB�Sꄨ>�e��ڦ���$��_��X�|��ez��a���u)%��|�qm3τ@�2פ�]F��?�W�J~x��諵/ۚ���4H�ה|�h*�ŗ�OyqI/6ۥ!�h��� A�̂����'V3���":ȍ���_����{�J$�+�"N�V�p�.6���5Op���ԣ�yR(��O�6��Lצ�᫢&�V�f����Ra�ڑcS�G�·�i6-:��M���V�|�Y����	J'�*Ȓ՟��l��1@��cd��WSHDK	x���l��T\%��=���7�ߴ22�̽��'�^�p�ź����D�iqw��|F=�H7k7�'�LW4�Һ��W���L!{�g!����
�JB=)��r6��Z4�vT���r��������X�\H� D[!o;��k������v�)��TdF,�AOJ5J�uscga!@� �Q���+��?��/��1��L������t�wI�g �g��gh�|�Bg���O�@��b��G��%u�1cXLT1���WgG�%GR��&N߳�X��N�h�Ҿ:�2 �.��$,*<�?���w������3{^#sm�igp*�ؑ
�Gu�����=ƾ85HT�mۯA}�ahT,����X�H�������uJQ׃�*Iތl��j����z��𷻿���?7M�bE^m&d��ib���^���{��Q��w��ax�1��C�&o׫~W9=����aoG9~~����jۖћw��䟴?�y"�X�o�����]5h��M�"��pU��<�H�#Oԇ0�G�N۷�ɬdGa�x,*;���3�65�;o�ċ乩9@SpðD��XyL�8���fO-{)sj_Z�� z�-�tQ0���c�+S�:��hP*g�0�N�2bm��u��Ŗ�)G7�����ن�@%��x��Gzi}�B��_����@1j��9yj&���ˊ�H51�[�8�͕ ���� ��Y�JHRx,�@@��3����(�ɰ�q_��PY�$�l/\)Yg~�$�~9������W�jo���P�QWcS�1�<�ʇ�
���Q�o%���cg�t��%���h^År_w��p��}?
�����Ե��ŕ]���V�A�?ޗ ��J��Y'ZW1��V[6v�)�"pܹ׳���M� �Pi�=`��<[���LzuV�o��x�"|��;%�f��"`�6U�C�
+(+�C��������>B"('�k?��R�GW��L�%;���?Q�1Q��}��	/��1����m���$=a�P�J���%�#����Kkd��Ï7r�vz����k����x�@�c��Ŀ���	����ը\+L��3���f��f�.��0 G��j�6�H�w��)��=#���&[N�QY575f��p/�� \��lv�`�2U؏<�ڕ�~��~��L;����5�ge�@o������f-�L�f�`7K��v���a8L;��P/�����=��3n^�PlGњjr�7D��[W#8C3}�'�[�w�k��'>[c�p�����=;W��^k�;u�2Z!b`�\�)����%輘�2��&n~��.��b���-o&d�1xHW[�͉��c���>��Z�o�W
�k'���<Ķ������q�˭̓�,�o�����.���\� ��of������R��dU�6���|��$�~Lt�A����Ir�i��P�-e�\muR�I��R�׏D�S�/p,L7@��C���Ҧ�y�Ѥ�h/SyܖV���
�o��Z���
1���wS�������,�2j��r��f� sz�!\�Ǥ`��y�$ƨ��u�xNQsNO힍a�*".�,���Wo>5^��>p�Ղ;�	A]��"���x�o"������$ks�������Wv��m��.'�K�˛��� �.�f���$u =�mzT���Xcbu��[�*�?|Hk
1e�ׯ�U	W��]	���8��G�ҏ�\&�Y'U�F��_��_�@v��zb�HY
���p�Ud��(A��'\�=
�H@�À���s@�*�d.9al峗���	�o2�6eQ(��FW��|%O�p8H�M�Ŧ�P%VI�э�\ȝ���*S>�fآ�s��7`f6�(M�A�#�8Л!6%,�$��[8 ��WMV�ys�n"����I cOco�����μ�o?(�<�}��A�1��"�R��
MH�ꀌ���+���ё*p3���<�+L���v�����]���#})h��ڜ�d\�c���A;���(�"�9�`LM�^��ʄ�#sZuZ��u��y�,_�������R^�`n^����W�k��Բ���WX���lq�5�D_��'�q�&�B��E��PSQ�ߗL?)����#ڈ#���[NB]׺	�8lO��`q�� �&8M�%T�٭�N2Y$_��Q���$��qJz�k�G�y�A��t=\��qƯK#����8�rh�|��+��'�'���G�7�w�}CJ��T哾���h�D�:	�pA,��_���Ss2��>Q��e�!��?�P�;�i�-�+G����t��z�1�1��T�Z/o�@H�C��0���9v��,pY��bx�X����*wt]¨�
���Fn~V�^�6LeV��RFIG�YDLn��,�I ңdF�'gG�߯5�Y� ,��/�~#�/SeN�Hy���w�t�[]n������S;0x���AmtUX�$a�a�-�UL#��7#�l.��c�d�:V�8~1~c�h�~jp:>e��n���<�Q:��Ǡ�I�H��yO^�٬R���Ί�YlW(�[4h�C�L��k�9E�tP�[��K�8�����Y�b��ĭj���x�I�&BD�u�� "� �i�*��/o��n[��-��-Ԓ���础c��`�K��B�G{Sȷ��}�L;{Q�%Ё�L�j��7騬C_3}�&�������ؓ��(��C����B2�(�ь��m!��e�G�E�h��g��*��Y&����[���
��Rn�Rށ�{
܊;�5�\9���|��RT&CI�����ٍ�f��][�����b���Ñc��X��ώh�2��A�>�����G0N��E�Ғ���v��8���8/��}i |����	�{�E9�)�s ��l'�mZ���rg���Gl�����N��-�w��4�92w/���{^u�÷9HU[:�.2Y�ч���B��j�Qu��%s��c���5ʒ��'	��ӝhh$��������Oz��q�$0�>��XbH݀�H�bY��*?_Q�,�J��^u�-3�?�Ǜz�$y+��|�5Z�����FѢ.B`2=B�+$�>�������jG���VB������Q�rB|{ë᪓�&�����F�˂�oS$��Y*�At�����	���2�¹���Y;���I�}��j��D�.�]M��^1��@\��j���h��K�Y�f�sC��t���E����mX�(�c?�܁�0!p|%� �~��ֿ���\��y��/hM,l��6�|�ǹ�@�֠����ҧ�R���uPC���W|J􍁡+
t�p~�����,�}�^^�բ���0�����8�C���&��9��yߝ�wf@�mv�,�&6�6H�����G8��@t}�n3j��I�����P`W@�Hdz`�M���c���h����`�9}(<@n��^��j�x�Y'σ���1�ljl`%U�b.�7�p��t��r~y
��C ��sP�wU���� &J��$B��ؙ&|5���ih��E�b��TV��;�0�3=-������:Ύ���`��<t��W�m�[zl��`r*�Ui(�$��a�̠8���`t�ݏÒ�0gވ��d+l��׽O=��x��G�P�ʐ�v��/���RM~�,'��N8�����mF��[M���I1_|ì��bk�
�nu����X��ef�O�j�7��~�9�ҁD 8������b���8����+v�|\.)P�r�]2R�<��Mr`iJwM*��3P+�r4&���	��#l����E��B����$\w�Ij���bٹ}s�rY:�6����:jy���[}�=@���z��8pZ��̩P4t*~��!����/ȣ5������+C�.~������P:{'ı�����/h>�	�MIBIƅ������l�io����E����S��h��S�C�@�D�U-u���њ��"bPq�ȭ�� �����ǡ����6�%��P3?��tf����� A@i� j��x%4�v3�u�3ٳ*��=�}���''�I�����v�L��0�=Ǝ�Ik3�T{�3��$�Yp[D���El.Z���]'��d���34���!�����(���?�%ZP4d�7�mRu�A{&i�|{�<�}�Ҕ�S�$W��l@
�/����
~���2�S�3O%)�{�1�o0�b���5/>N.&��3���~��b��*[�F1˴Y/�^ߋvԐC�V�g�/x�Áz]k<2���UƴfaO��³xI�<3���'*$�bM���r7A( �������ݦrZ��q��W�y'Qٲ�1/�Y#��K�I�O�kˈ��N%Ƥ�6ھ7pP���>��wU(=�f*�S�-A�L����\�v��cC6�C֫�*/��@�A_9�uat-���6��.\�ʬ��0�sbq�]�Q,�|�%G��\>*
���v�ƍ�O�~j����~�K�����[��U�!�Ag�*�
�l-s���kTh��/��1�;�Ϗ,��<��v�S��w�١�����������,�޸ ������������9�|��?�83f\���e�?Շ� ���Lv��,^"�J&�guk!��	`S4�%>R�����D%�Ŵb�_��hJ�$+��%�#Wq���S͘�1:i�,�ͪdlll�Q���5	���\�w�Ks_��W<�u�Ɛ83ƚ���n�b��B��&'O�o�}�8��iڮ�f���:dB�kg�~��[�?��:IW8�ֶA�7�����=��)a�K�h��8��@�x�&Ǣ���m5yc[��T**ۆ'L�9��Yn���'jz�:dD�a��$�\���T�&�Ba8�	;������Z ����>���MW<�ڮ�簻N�`�ků3�����`i�ۨ/�ϩ��G�kw٢J+�C��z![�T������hR����C�H����K����/��l¦+#��-��tw|���,e�xK�\��G�`!�$�$�R� D2�mk������Z��ip)p�p9�<0��	�h�SSN* ]) Q���2Z�-[��h���b��r���:�c�3���c�3�/�����S/��X(	P:,��n�V*��Z�r�t�Gkj�j'$���LX��痶�4�o3���"ё�?R��� 9ɋ�u��ͧ� �ed[<��̔%`y`�a�F+�
6�����F��46�x�W��j0\ }�yy��˂/Q�¦��rA	�}��4�6@�Pa�^6!sHЩ���8+��?�����*��ĊT���]��켥�$�0�X�4�Gc=7�x���8����@�00��\cx���>���P}�tp����J��P}�4���pv�M� �K�a�
t�#�V�de��S�LI����iǢ5(W�V�Rm:���1v���_H��)�>MNC�ʏ2�{Ŏ�������C�q�I�������6���" C'?
��K0"�0���`�j袇�b��%�P���ek����2h�����rB���,�Q4B���l���\& TV��_���.ÎHek��]l����<����������^	�G1{�.]�����բb��a�7�.�2���iC���n5�pu�V��ݚi��/������a��JK�?5��2�j���"O{��6oU���l�R�f=!j�Z��tm}���)ϭ�����%m'�ɘ3�"��P��Q���B���y����w�B����� �Ir�nw�"��U�,�#^�(�p�HP��#贮�]�#���8���3/zc�_-2p�)�ɹP����jj��������]���PZ��Mp\Ρ��yQ����'_�P����Xl�to���r�`8�sA��,��������ϒp/8����'*&y��c����9��U<��l���x������g�qv���cw�tX������B"�yq��/#��UEjꂧ֍>�-A�v�4W��7�×&'p����&~1k!PR�?|N�cp*�zPΊe�1�Z��;���8̹VNP�g��8~�~�",��q1���7�Fo�z���p0�]�^S�B�a�o���н��ʖ����~S�T���`���+-�를�8ˌ�\���P?�t�����<ZY�ig�P��j�W�؉A��Д�ј���ET�c�U�wD?C�>2x}�	�����8w;³38i�!��Ԯ|�HElP����b7�(O+��n����n�ۊ����5��v%��h�F,JƓs2��Z ���~LY�aD�~V��ӷ�[W19�@qk������ٹ�6��n���V+5,��l4v{й�Y�y#Ʊ�w��ۢ��Z�^d�9�B�7ü���d�!
��т�Y�r2K��W�񓏢Vi}��Tɬ�\��0l:#f�����h�T����1����/.�oA���=V j�[����:��_$���ml��-�(�lFKփ��Dٔ6��{Xsn{Uch�	�X�+���ۍ7��3M�Y5j�aI�<2�r`
�`�iYȻ�,�,���e��B����Z����*p����1IP�]���ш"c��K�&ڻ�Ԗ��D|7���eC+�r�:������<��9ԓ��W��z�����]puA��r��J���oe߶!t�(��]�dDk<+���\\�8	QAѵ��,��/2V�� @�x����C�<�Z�S^���π[$��Kn�m��+�5�d{�����)�-��1���A�Ԁ?�Zܲ��0Q�k��v8a�����=4�� y� ��)&��t3�]�2��5��^��6�0��W�b�h�u��#[�e�E �=�SVcB�3���M�����w�
���
Z�_����k �&Y�/�k��n��Оb� ZU*M��=MK҉�G�rd��Y�m�n����
�i�	���~�8��������%N����uky�R92�C3���?�d��w�`���}�?��=<�|�:�5��j�jɌ�Q�ؑ�9$��G�����uO����m^P�t���c��|/��5 �|���93oE2[�`E���|�����~\��o��F4H�/cb�˲�W���W�b �y�koOg��p_ �����m�+HƬ�E�|]�HЧ�E�F8���O�f���eI�3��^�0g&l���9��G�/��	�A��6��eJ�]A���n�Y���;}��K��t���Ӡ�c�^$�-T��W-.�]/m�����$�9�d�_V�l[}e#�9���G������%65�0��(^�+���B&�}	��%��G�1��Y���̛��0�FP=��7�:D�H��k����
F�z�1��4Y�LD2�h�D���yRfG\! ������.A�;0��f!�^NUz�PL��2��7L�n�i#�o(��)����,�Hw�\+��Zm!Nt�M��5��86�:�)�fd��&����%:ǜt�6�R&�[	Ѻt��q"h�jQ �l�-�$��.i���EL����j��gޑ���ݏZe��X��~�o��dz��6zAQ��v00�c������YMU�z�P�Q��v*�y
�'��p�����j�*���`$U,}��z9��t��I�תL@]x� 6W�̘«L�������0]vs�ED��Q p�6/�I�Hx������ S���
��������� ��SĔ���2�H�����J���cÃ�3�EHғ?_yf�wɍV)����f���a�nE�"�Y��<䑫��D��j"�@8�5�)�l��J		Jh���(�B�GZ���B��P�ٸۿ�M��������0���FC8���{��`}��� 9YȚ��^�|g=�>%��ioǙ�% ��u���@�?��Z�ր4f�(�Bx���:�]��M�e2#��d7Y����C���ynҚP<���kA�����@��������_�t��x��� �xww:r4"*�y�T��Ѣ2�D+��F9K�Ĉ�
�D�ck�A���QG�&
a��br���b+�{�{J:�����w��E5E:V�A�^ڒ�Z�!�L��w�|L��N�����-SV�pK��w��u��j�^�31G�j�ze_WlR�&V(͞�oX��;w�AGB�շS�f�y!,1h�u0�5II(|i���4OϠ"�p�K��g�%^�!��Cu(W g��!��Dݳ���J���gZE��Pǵ�3�[�(>�)KӴ�R��R�G��.;�Oy�>�<���O��R iD�(6������F�fx:�(�!x���8���ӥ;�:PP��&���3�ՙ}O^]�Ţϥ�Pw�ͪ|僮�C㘃_�]�$�bH��P��Z�`�HK��=i�`3��m^q-�3J́Hq>��[��Q�1h��+�]�e���P���&��w#;j͇�h�V�g,��7 4���~����� ��@gp��Ze/�K!ӕ��mt')��Xb&'���F%�H����: y#A�FuH$��_2b&���h����?Yg���A�c��m#h�) x��z�wJk���6����yQ��a����r /D��ϓīiU��_܆��e��)��~��-���mD��⯽��d6�u��yֆ���\�R�q�T����Sn��@C����(�7�rʔ��O�zƝ$O���3zL�QHv�h���Fy��o���	��ZY�Y`� �e��#��}�ﲥ��`e	'W��^��ぞ����t&�%2޹�E"!Ot 'S�H����=?*[���(����tn�B�Q�y{ӝoW�{ch��A��¯\��x�Ա�K��>9����e��Bb��I���I���"B�Y$Eā[!p��o���+�u���د�'[ 翵�<yADq`שڪSh���;k������5�d�o��,�^}0�,�x�{0�6��d��5Ӡ�|�Ȝ-��.c	���l6_�A<7R�b�S�-�tp��pM5�){[ŌE�/���5_Nq�.����p-�K��H���׉/	j�5�甆���Ź	�����xۜ{�e�����{�?�x��^P���4���e�FΜAwn�x(D!!�F꿍
�jH{�Hs�ac�d��h9TS��&`��u����4)ݤ�k~�Ǻ�!�-C��E�-`tJZ�Y��t�ȭ�#���k|~�Ԥ� 3�0)��Ov�����:���揿S�Ʒ ���+�#�B��z�P7�T�nbZ+�{�B�Л�d�ri�0�� ���K?g"� �(��
B^]�Fj��%[ܳ> a�}Q��$�k�'�c��f����ǆB�I���J���%QUԝ7����	��@x�_��d��ȋL���.�ö,nX{�[� ��8`�j�[�v���֨S��]]NI�����wYN7-5�Rd�ho<��\�JK��4�0M���:]2���;[�C����_�u��� !3N�7�����u�FAPq��/J�h���\�
:}�9���2(�lx����KЧ�j�� �9h�w)�J��7���)��`�qL�]=�e����.9���ԅ
k�L*���Z`�ߧj�PH'�Cʢ��(VX� r^���
ji-��]"�����820�І���E�t���Sq4nRm�buĀ?mFet����Z�T�l���̬y;��E�-%�*�
RO�ӽ�܆�+ݘ�;�/θ�oU���g�)�L�_0�wH�8��Lޟ�&5��$�
"z�>��q�n��F�7Ψ��$��I�o�B� �4�"?~�l6k�N���RUٿ���%ڠ�<1�P���N�p2��Є$ПMY�c5�KH%�����#	�s���J�a J~9>�*G�d�aB
 �1�c�j�<D�b*^�J�4g��Fو��h#(T�?>��	�&+�Uk�V܉� ��'���L�3���1�$��9�W#s1���,�x��&�����mHWcpʋ��*����>�fM��[�&��ё=��u�m`O�\|�.e�� ��a�-��O߮��ߏٓ��/g`i�a�*�-Ci�6J-8���^R;D���OR�hFQ�����P����=1_(�ʸ���˳��,��r�}R���H� a%���凒��Hz���~�jyR���������M�˨��{+}h���	Q�������[��6��O�W���g�hi���}�;2��U*��?(����=�`� g&_�x�6�l�^n�h�[R*�7%.W��>0l��,E���j�V������l�*KA��Fx^,-L��ϏbK\�-��zG���I�S��*�o�8�uKTg�("���c2W�<��sb��o��0��z�u&�g+4�۴u�Μ6���X-y|Ε�0j�]�+���9c�|Zq�*�-�Ώ{�k �ᦵ��ܫ[�Q������ �3� ����U`~7�c'�/�UU���qӷ���u9�}"٧H�>��4��Xf-��eՓ��2�롛�x��@Ho�$:�����<��膔��j��n��~D��y@_��SG���d�N������[xo��I�.��X���k$�ڡ�J&i	b�������|�h.c�x#�و�����TL=n x��D��q�sOR��nI���w^�a��+�E�=��=�����(SG4)\�O���nT2��w����wA6J��}�RdF��P;�ǭY��\�GHG[;���4�U��_Z_�= x��ێ˹ ���w������%#��7Éx�`3 �:j�������
Wus�/��T��7J�@�=����7�o�[6T}�h4�����[E����G�a<����!��1pg�@��K�R�K��1�l��-��xȁ�龐�,25�XŰ>^���c�m�g�i�$�Izu�c3�̕���H�L�SB���uhyZ����Q�,1nuTܸ��m�R㤸��XV�$�ݨ��'���Wt���P�&����� ���W�2�{gf�C��W�C<¾?��^v�_O}��%��_)@��7�H���G-`Z��h�jr-8�ڸ��<m�5�e�Qy��^I���/�* A77:�v;��k��0�D��(�vkH2�}p���2�j����W�?M�mq������X�ƤR�Θ5��(1��i�ሣk�����eu�!�'�)�$<'�f�Y�z������5f�����$?|iv0!�wJ�Q! ��8��� ?i��۪4`8�g��R����V$C�}��cwW���%�=��dk)=�#k��½+?�f������Z�g�6�� G`��UA���j�Hg�=9gx*���}i���X��}���"% �D�1�]hܪ�t��C�vLw����<����3RSA�!�a��"E%:UB�\lG�쿝9�W��Q{�'_;�1���B�n����CY�D}r��Ȑֱgˁd�Xʓ��6nCGE�!؂M�ї��{.T]B>1r�GmDX��$�ʸ������R��������"-��X��+1d��]c���\�V�eh�w#�����yv����A��a@��bѤ�V��7�h��wqM�A���[ԯ89�)Mլn ��Y�#��i�3O�-��H�O�#��'\ƼB}��LB��	R��]Ui8���۶xv1��|ƩF��:p �+7�H.�"m��x��.���/���$.�����(H/�0X�5�+L*H���k��=�<�so�������Y%�3'�p�2R\b��q�Zࢁm<9��M�
F����&0���2��-��g���y���v��s��?�^ ������=4����WHj J��9�E�[�9��C��M�6
F~F/ە$aa5���*�Rt�tFP��W꾘�-e�(�-!@�G�%��-���s](��0��Ld�ޚ�Ц�mjm}� 9:H:n\d�eAux��Ǹ��t=� �o�����1�&��L@�^ R��3e��%տ���1�(�x&����ySp��]��86���T�V��H�5�qca�X�6�Q�k���rEW;:�^5 �ޙdF��tF&Y��FY�݃c�p�gt*�Lܪ$=m�m�>��9�۰����qS+2���d1�b�\��.��z�ܛ�<�~*T\�L\\^�:Q!C��<O�_��e[ɞaQ��\"WKfQ��2��ƑP�k��x�*�"��BJs;�橛��q�OSN_��a�T$ܭ�5�F��Y�e���,z#��0��t�Q�×��}�l�v��a8��)�6 ���u�ؽ5R�0�Np�E05q�i>P�鳕��kJ�]|Oo��݌Q��x.V�X�9*�٠�Q-��Y��ٰ
e��O�Eڌ��63H6Ld65���g(�pί��@�K c�y3�Ȇ_�Ù��Јl<g�m��L����\��I��&���rq�a_�9�X�4D��04�u�8N�=�G�P%�+$��_f7kn����Pv�us��Y4`$���(k�T	aV�Ӝ����B����);b��A��ؒ9�cz�5�u	��'����>_��O?�2�+�7��Ů%~C\�j��4���ot�\?�s��ۈ��:?rZ8�odM�&��`I�T�r6צ����ъ݌Q�!geӎS��5�d�jv�&���JUvJP����C?���s��n?`�T���߻��t	�W&VՎ]@�d�]ӱW���-t�]��%�ҍ�sVP@�����1-	3A���7���O�ߋu+ )����L�����IDo$Z�垢;�0D��kgۖb&d���[8�8��a��~UZ`3E��)��6J%�9�"N;���Ȗ~�%u��|�6��T'��_R;�0I]�����˪'XRbl�%�{�MZ�>� t����z+x�5��dA	���6 $����W�y��g�/��9gU5����y/K�h��KIo�')�mӤ!��*������������d��ɴ+��v�q�姸�o�*t�?�b�A9��YK�	cM�W�&��J
l
�s�y�2�n`�L��c�)N���sQ���ut��|���q��}�]#Bd�HXB��n���A�I�4����Y܆�-���W����^Љx�L6 kߜr��OF��_C>��J�	�)�W}%�;��0��������%��(�X1�.Uj��y>̐�ql��QT��l�_��h?D�n7�zJP��cL|.�q�u�V��q��l���#w�Ԃ�@�i�z@hAD�*�,ԧ5F�qT�"Ѩ2o���r%y<��0�"(X-^�{1�(��!t��E�v�1�K�V5��P����K�&|*CN{q`��i#���}���{s�W7���_���>~��? ��n���U<���ľj�Π�6�����2�m�L�%N��II�`��=��nCI�?+� mԜ�V6jte����<�:y�R�;���>|B(U��n��튧�!B���<C�.��r:�RN���A�)���ڐ�,���S�g��+�
�P:�{��� ��;�`E䠴 vϤ/�ls�,Kk��?{Y�T���U�`!E�=�g�²/�v�;���t�N� -(c�h�te�p?�i;�[��9w)Z�O@PӼ<�^����r�B����!S�8w$y����XD.�R������:�\�o��%*��B���r�J"	rq�P�!B'�]�·�=1�/=�+����bh���pb-��x��P.���#"���|y�F��k�^��je�8P�Xi̪�))������>N�	t�%��ʹ���%���xN�xC�]$
�a�g2k�����ϐ��0���7{���h�_fŧ;��V�Ӣ��]x��Y}��MMB�%(AEm+���'��#A_��K�������O�b$IZ�3���h�7l0Z�� �f�WGz������(�O�ڡndhT�v�vB递�*�����V�ϦB-����A���c ^S1q�K�]�F"���ꮦ���9�z*Ӆ�����I���;�nNQQk+U�yV�����\�KxnvI`���
;ϟd���ku���%|zR�0�I�U"��{��W�+>�r����J��%�l<���C3�) �"��(�iX9z�f]vU����=\�3`�Y�28���1�j���Cǡ�vӨQ'�Cb�����[���аҫ��YKf*3���r����2�m��k�s�=tq�|���R�Í��m>�;�e�us5��J٩B�)ə�����qɢ;���lq�A}����=6��O��'惴�m:����!x���̭]�|Zv�w�r 5U�i�(�5����1��r?v�p���&ìW?���/��~���"���qz<QB�D�,;y�j{��?+�g������;�(,�i�3[�j�J��kW��٭�~��:9tt��b�Ƃ5>���b]��3���'Y�}Nf[���͛ ?����j�h�L��%H�F��Q�Vm�����q�u�N<+1#��F���զ�m���hb=�1�"�Yr2?
M�R��\��e��i|X:�h�͍�T�2e`�`�9�_��)��i�*n��^�aD�
�C�ž���K0��1�g���Ӆ�V&ӷ��S�RrsP:E���>�u.��(gq��vSS{A�`iZ�VX�l��0]�j.-���HT��փ�8ኘ�e�	8�Ff�H�#���{2cO'>A]���ɐr��G�{g;�� �[��L�e҄_�>�j�&�"��ذ�����&��\�`�
i5�:t)�hZց`$�3n��=���
�2B<9a�M�R�8�~��A����ڕ�spB��q�㷉��vB�|?�
�&4�:ԅL)��{t�]�pNmt�� ϡ��k��{6}h���셵�{b�@���b�⯸����-���Ǝ�������V����<ǝ�'��2~hߗ�f����+�LEL�C��y�_�5��w�Q�5Y�����8�O~r2�a��>M��	����3 au��/i��XzPv���x���?>�y�)&��f�>v��լa�^����M�碮��d�ա�� ���Lg(��Z�P;t��x*�aP�/�[!MsnA$�̝~Ws{�t/%h�˯�>0�-Bl{�׻��������N�q��'ɭ��@�"4�P5�>@b����77	�/�����ؠ��/�G=���HEjR���"�1����i�����_F�˛6�I<��M]���Bۧ{���C��˵��r�A����Ʋ^����l�ڏ��n��ke�gI�a��ñ�+E�)+�o�<���^���*'$:3��5�K1��_��S�r.k�k�[5����Xe@mO��@&%L�;M3P�J�����C?�;��v��X|c�$c��_OE}B���[pnx�T���*{�g*�sGO%"�zR�w��ɘ��C��
)������+�#J��h���Lij}�{�,A�,< �uO�c(�D���f�q�9�׮D:z�Ygtw��馭���w�mz�@�b�4�ފ�Un�h�M�l^�F;��Z��ދcJ�nՊioA�ۗ^p5f� <�}��9;�1F����UP931�氟�SÃ��`2M���MI�9,8T	�(�����+����ZP5����bQu�R���#�W7�=.�4A���CAB
q��1�_��|� ��_"��,����I~Z���	eO�~;�M��,/~r�d������3#;�N}�Z����+�3��J���N�d��F�w�sK���R����3���z�үْ96r�䬗^O7jƳ7�|D�/Y��Ǝ{�{�IVEH��wS�xg_��M*9i�B�s8���q%qW�� �V�$��]Y��8�*�����Ǜ�~�'��^��]���k\�#۫˩8ܵ��kZ$_r�;`K݄�:1�˒���W�R�I�&��R2�{���1�zuo+BI=�Y}���4�W�#���׵��,��P�4�?�Z����A��%�'�w��Cz��\!t]r��1��*�Gu�x�.R)k_Y��a=㤽��O���?����*J�pX��Y���7x��?�)�� ��fK1�h�J����lY��V3[�b��TU%(�~�'�20L8T��9v�L�[>���{��҃���p$֗�j+UF8�ҝL)2��EA����}���֘����0@���=���|���$�r��>n��}Sr ���AA0M,}���Ř������7w�-u3Wa�tkVV�(����I�t��4�熄 ~�0r'�*��\f�l��1G����������>qo%)%�r���q�o�+9h�Z.����V�7���>�
���?R�C�<�4�.���k�V�n
:��fy��m�P�#���V�jva}��e�w�w1U-�$�:s��NOl�gX!�,����*�|%v'\��T��L5�@�֌���C���&&��Jw��*�pZ�����e|t�p�� ��:�nS�a�-m�@��J��m���$<eV�ίHYa�*��uK;"���EamV�.~'w�����G�	
7���hZ�B�o���ș�eC)��Jk����0P`)��<���V^M�GC��
��"�3"/��|�>�?����'b|dٟb�[���N/�U��p̮J�$n�$���-1ꡫ��/t5!�\�F�$k}f���#F�7���Ҳ�v��&���r��%jH}79{�[�4����HH@j2���h���Y�?�7�M]4��wA�H�: ��@:{~i���`r����4�bT�e`o�DC@�?'���a�1�F'��)g�d6pPO�u'I�[�S�\����		�{)Bw��	��l�#}�o?pĹ��h��Q����~���c��**����F{�UM�n�w���V,�QS��I|G�%��,����m�Ȩ˗8��g�dgI"R����x�A�-����1ouܙ��r�s����nX�+��)`
;dXl��k�j�u����r&���G慁;j�E4|W��g���4�aA�-�D.�tE���f�3�:gtUC�>�^�W�\�=��릫Go��.��X��T=hR.s	'�pUH��ޭzKD�� ���p��f��7�o:��S;����è�&�פ���ݫ��N��gI�Ʌ{Q�k4D���9i�4c�v��H���8����FVC�����I	�8<(�5���auA���QOI���k%��'*,�#�:�c%��6ѐx��ȀF3��p�O�</�0��Tp���lg�d����>�"��knh�x����Wr��W1�Ƶ,P�1GT����4��(�3��q��Oq����o�:�N%��|̐c��)�s���^�6��u�!<���P'���c�ۭo�}C^�z,z_���v[+�^�D���P�{ǅߣ�v)�{��l��E���(�/�]���X���:���)s��r�8��]�9�aֳ����P ~+��CS��ӧ����	�O���$�]l="���g*b8�Y�����6��g;�~�l]�:8,zN���>GRAL���$}�u��m��t���y�$�Iܮ������&i�������/��v��n��^�2��L*pV��Ä�"�y�(2U�E��*�L���hF>9� 0�S��@#ƥ�z�yIK�p�g{���1T�J��E�\���:�<�՞��st�a5~c�Z��Y.�[�
B�4�ge<�#��F�i!���V������D{؃�v�ũZ���]�n�i.rd,R;�)�f�/��Sy5-�8������~PQ�z�ٯ��������9������5�Q1 S`���8:��ʘ�W�g�D�.�����S(#`% ��9\Ǽ�{�Ox_���%�%n�UI����T₍P�Aڲچ͂��K��ꗘ��-�ӥA�� ��]�c`��(��'����k��Q6�{���$98N��xÞ-y�e}��a��T^��:�������HW�B0K�\������zJ�i4�Z}����@_�Wzw�@p�!��H:��$OB(u�"ӌO��˰��I[�"l��B	C�W��@�s8[V�;(rԷ�A�؈*:B)zIiG (��;��a|��C���:��(�<_�a�m.+P�ѓ�Ɂ�p�&k
e����PMUq���]��8��c��!�XD���h�9�f�3rf���8%ʹ�08�dF��l^�	5�~S�����8�΃��|;��%��:��4*�)J������8�ɧ�r��(
�^Q�O��%��I���������\WK�K��c�yV!6D�-@ÿ�j�*��j��x�D}���f{�/d���� ٠j�\�')^�wv?]���>�C^��͋����wη�C��#=8ص܏,x=��ç=�{v�S���梠/ö=�U�eTDT��ey%��s�Z�0$�-@Ņ,�j��Q�9:�+���ڇ�ά���G,n�Ƣo|;�tWˤ������� �w�k[ȫrs���xM*��ס]9e��7�n7��̨c@N�5��A�񇐛Y�$7�v+Lo��rG�ՙǙ�a�቏cp?��������r �H���E���l�5���Qe'hZ�pj���ls�2�t�%-�dK I�xP��4 �`��0�����Q�k� ��B.ۆ���!\μ]�B�4u����\���2L�8�2�a�D�<I j��HtW���<*ʱ��8�td��j~±�]+�H������V*i��‑QwYx�p���^�Ө�(�d@[.�T8 �p�9�SM� �轉�H��c������������.y��0}���&�UT��ՉT�P���,}��AH�&!9�zk�?�>g$�X�mOl��� ���\d��2��3�=�� �+#�2�/pv$ �(>��o)_9/߷�j��|Щ�����	7��qԚr N�OOD��V-�)*���9��ʌ��¦��զ�-�d�@�Ji����[o35�e�Q�����r����I���N��&�˖7�~�e��V8j�v���$݊��@u@�o���֟����4a�����N�#���C���*��vj�mK|�0O���@���l�[����)�}0n���f��y��ߟJ; �=��4-<�?.����b��j��y�!���qF�#����.�C|4s,q�����݀�$��)C���يMڣ� ��MP��׹\*"���M�+������gxW�x�4BW�϶7$��P}��'�lv�8�P�aS�+����d�3M�7~��u�g7c�,O���X}�Ҿ�5�.�QNH�k{��i(�~(�9%(�q��� ��,%ϓ����c�8#��ԤQ={
-��`>,8���_s��8Җ��V)o-��NȂi#y:5|G��H.��R��s�0�ޟ<�'��M��'�sy&3n�l��;����Ic�t�d�J�on`��Lgn�k8F�Z���F�B��K���}}�r�#�d���ݠ��B��@[9���:+�5S�Pba܌XL�=����s���9g��\�~����&Wن����8��z��aB�Te��P��0�(�G��[�ڜjG��t�b^L�If���z���j=�~���6����1oW�7��5r?��ú�>>��b�l�?��,��Xĩt
-6y2K�`�Xv6VS��.S��`����:Au±!�*8�҈.�ۏh�����!m�XyG\n�����k��13�������>^�q���vC
;m8:���}ז]��H3�b�>�[&�Zeç0�C%B���̭�	������8z�������^z�%f$�po%:��f3��-�,#�713�C��QC�X���12������"榽w�$����#m�1��e��J�OJ8^�V-��I�j�S�	��.���k���@�Vio'~!P�n�A������-��~v��qGӳO<�XU̦� �9� ��%�1`����g1{(硿?�O����mp����k�U���;��YЮԣ���(Ƙѕ�E���hY�<�da:$�}ä���( >^$"�� B$�n�]�}�<P�	4P(��m��g�_|,���S��.Ex_Bv�����vq��đ�!'�PJG���ݵ�b
z��]�W���u� �����#�Bc�J�.���Mn��I�2�>�S��G_F��
k��"����M�ǝH��/MD^(�n���T����q���#D:s4j�ئI6�G]��/
��΂�:�&Z�߂P9�ʦ�7H909�5�[�ז[ ^h�@���ew��r��ȃ�ڍp� ���g���	"�G��J���9���^���)�T��;F~����C�=���u�#�~�O���$bl�N%�$@ �������`��
p�d�U1�U��s6*r7�֖(�~����p���KG����+Ɯ��5j���D�7�Do�{q^8O��$K��~^9&O��+�Q��(g��5������'}@�)�ȵ:��Y?�g{���M�zF����`�&j����{��(���7~�'s
\֠;o6�Y�#C��_�v���4v�}Ci�eQ�����W75�����������CBm=������-x;�b����K�U�*:SU���J� q�����*W��t��v#�4x�Rx����&_ �-B�Y2r��Ki�bw�����2��߅f��c�a|�[�t��=����\I�!Ѝ���������{Bf����T$�%�7$L��  �
�W�mȞPCU�#w�R��BN�1 =�ٳ<�<���f��UO7
�������!rhSc��X���`���ʩ����!�$\�'��q��DU�H��q�� %ʫ)�D.�Y3�%�$�A�A���et&�c���~ W�d�s,a7�֔��?񷷀y�0qU'nS���HM}�g�Ԃ�i���K�j�!+aiȘ��$D?п۰�qZA/e{������L����7y�����{ʌ��CS1�q�dw��'.ޤ'U��Յ̞�j_ �%F����ڹE�UO����\������ �°�\�U����nfjw�xx(��jß�L�,���j�l������n������;޺�%Ά��;�vL~�RK��/(�s���7m���O�F�ř*S��@4�R��F�َ��4Rx���F>#���f��	H���\-�������V���|>D ��(� 9�N����,��R�L�=�����߾�<ƅ���O:�_)�����g<�Nծ�P�2?݌�E�u�d��m�Γ�������P$�� �j�bb��v�#��*+����q2��Dl<⃊U��qY�D'�U,�,�6��j���v�Υg��I_�7���&{� �BG��A{ծle�-�-��O謒���-�h�}�Y�֘�؆�����;�j1y"�7�EB�i�x/96�ѿZ�?���i���P�����W����� ��%_�@�XL�d��_[�/{����f-��_�N�L�UROA�NA}��tфW��Z� /g�T|��o�۵���H�ԯ�#z�h+Q���+X�⨕�l¶�3��$.�4̫y���p��㠖g1����7Yg�F''O�'Kă�O�gV��K�'9�ȏM@*hT���]4|zd�o�*%^�5ѧ�ǒ��T>A��f^�"���Z	Z���n��+�;�Q�|���@4�ֿz�@��XP&[�Q����"�j_M�g����Y,�z�ڼ��%��Eg�9�q>{iQZ[��C����<�g���Y_�gM�`7�&6��w^���QV�MT��F�ҏ��.��/�B���jH`#�#$�sg\ɷ۾2x>z6�u�L���#eo��9ce�ͯ��@���\��υ#@YgLU���"Q�/㛾(���307��	�m��/�My:6Kh��:�M���*�~.2�Bf��Oݻ�
 M:lɺd��AEZn���$�~X��坃;���S��_l�i�������6����?��\����~a`��d���L�3�{�� ���*g?�\I�p�!�ꦘ��K�i��P���t�����̩x
��W����EtE��]P����C@����V��'Djŀ��,fw���2Y��1ǹ��4�C.��P�~�J���5.��w4��vR<E:��BXO��A,�>�h桨=#�_`
����ׅ�9�������!�YI�2��wXE0)+�M� �W�'&.��_r�t0�4|�x�J��~��e�HD���k��y�	��a�=�]�8��C6��.�p&�4�`��.����{������3>�^[v�2�"�g�(�+¬�;�CԚ
^	�T�!%a�����[1�9C~�=r�Hnk�D�Sq�<�o�r7�h�Ϊ����E��u�&���P?�%\���f������{�ߗ8 �Z@�g�����+ό��=����Iv�f�I��ұr���������~w�#<--��� '�OEwi��\�1-��<����?�I4�l���?h����>ܹ�~�J����Kk�	@d?�.'Pi4�R�����˫�T>8������N\"2*�y+q��a��o��%}�&��C�5_�6z)��x����W��j� u��r�2A���lpW���d�Y	mY���י���7	��p��Q�GM<��q� 2�!:��|[���k�e��uYe�p�W�y���e1{�?��
�U���>x� �0����RSrY��Q$�^Zu�e��������.4�*�i-��J@��O�w�:�L�c�.�эM`�ײ����:��w���㒾��Wg�׭S ��)��?KE���@2 �?� @s=�I�f8�:�d���f�}��(�ӥy��m��=��`G��0u#��cR��-��/%�j�x�����$�ӡ���j����F��9�Q��	���q��EZ �x�;Tw��;L��sѷ��֡�k*�	5ڏ�!��vxXo��ߟ�\	��ک�s��q�Q[���O�T�Ju�q~���j�X���)�jd�5]x � �@"(w$�P�'BT��� VJm~M �Œ<���Y�.@2��x~���K��	,^�X`��Zh75JI(�'�]X���?�H�
��gܱp�R�Б��3���r�#,�� /���ȣ�^���l��/8=ʡw>r8^���C95|��)�8;���l�bk<J��-�>C�.����,�)���&�%�%k�>���xﳭ��� Wp�sv�����@Cf�e��' &�x���W�����uk�-�����~ \!o�ZJZ��[�eF�|�vzo�֍��B��EX+>���J`��̔[�<qn&_�w}uo�F�$58�������(��;}�Ӆ��kg�c�>�����"�������Xt��E�[�w�]
��(?C�L�N�̙���W� H������Cl�Ht$���� Z���WD�Y�%�</��8>r-h�|���-3_�Q���B�	���C�6}QX��S��gH�a���(�xn�f�l�.�
.s��Z�����c�7�al��N�~���0��ub�F8��;���@��	�cnT]����պ�73.�]K7��ZB�X�s�k�����}��Bu�v�lZtݼ��|���[��lX��"�
�chB�V�(����*�fC��j�6_���){th���_�4���C�$����d/m&W%�r�F, l�Hc�?�L� ��St::{ D��m��@p]G��Pک�	���=����q�l�S_q$˱����﹙.+��1O6\�*�umAω�Q6Y�;L�cW���fDx�0�-?q��4b-s�w�9�<ث�T}V��M4�8�G�V�n�h� e�1�N����9�f�ɑƀ���eNJ���{I9C�~�|}����rۚ7k�=��`���*�j�oOgQ�&�s�t�YX��~�@��2{��4�Hr��7���/O�2,���P<C����r Q��φ�Yf�O{���ޚ��~@G��B�*BDR>L��/����$�����@9TG��,r�OU��������-���m���YM�c�ԢsI��3�@���-g�9�-cE \���Rl�����_���J�QuJ��[�m��C�;��>��"�*���R��a>fgۻ~UU��1���ϊ��6��h�����*�-��D�)Sa�t�"���ϥ�S0�߾M&�"�Z[AIM�rR�"��o(·�MG,���-��nNՌS��8_�2�.CI�QAt����+�\3��b)Bω/Y���H����Ong�8�1-�LJ��?�Op��ĨU�~s��^m�#^PP��M.&a��=,��3���fh��^i ���܏a����y��а�ږm4�*��L�`ij,KS.R��N'��D�cuV`T���>r:D�gP�	����Äz�Q�pE�!�p
�ANd��c�5��8��T��$��ɇ?�5�t��|�����#ɮ�-7T�3��
Ɍ�V��d25'lߨ�0���5��\	/$.�K�7�Ba��Ma��"e������Ǎz��@>@���i���ܘ�F�v�CIQ���h��,U�����lg��Oo_=�����
[�~��T��1�im�>W+�eyq壸��Adse�Phsں�AMF*����f��`t�������7�T��*J~�4��]e��7?L:�_1j����K�n쟪v0�/�Ǳ���QB<d��d���XVMn٩��}|)̇�1}S��1�)PO�ל��Z����Rҳ�׍�	B*�O8#�|b��#�]uX�E��� �e�IzNK�/}��si`�:��Y��i)��SMhP�
W.�;2�΀a��R��%����j؆L{c9�6_g{��I�Ǣ��*x�Я.X%���	��&��kl�F)AN�4�,�S
��'��$ˋ�m���n���I��d�=��[N�d�~P�?�՝�nQ)ZH6'(>R�8<���2*��`��= ���2��"@���pf@��^f��3	�>�����������;��т�떁9��Cn�k�a��lg�E۫: �➹j��'?+�}��L��Pݑ*�$�+x�r�2��i(���ʻ4���	�fQ�y~�	EZaq	iC��0jhk�*@u�#	�?uN��Kf�m�k<Ϣ=��ȇ�����$�\�7��1�gs��	���c��y����nݍ��d%���|�����h�\nm����Ʉ��/����y8����4#?(�3;4	?N�W�1w�����_gd9�2;���Q��A��t��Kf�A��nwMh�N�:n�Z��gG���剨\��I�ʃ���C�=;�k�U���FnL���n��l��R���U麍m�3e\�[�����x��;�JK�\�=���@j?������w�sP�œ�C��W'��S��F��M�G�I鏓Q,N�@֥��#]����t�C ]�F�P����8Ǽ-:D�Z��x	Z�Y�\C�!e�y\�ڵ�Y�F���O�m�vh�n�f� G��­���}��m87Ud�c��3H��=�����ў�x�#v7�SG�sX���)�Q��h/E�S��2zjM�� ��jB50����Rg�$�2��;f�/=\�����L�K! �����e=P�4"��F�v��MJ(���NV�V{Y5/��J�NڿB�G:�4>�д�%	�&��$W"( ��u�XG=��³��5}M��mˤ�z���U*��[;��|K���]�����՟�%���LH�`5죏Ǩ'W��E�Q�vA|�#�[Y�*�����;��]C���Z6�ه�G�ISen Vei)]�v�l�c�ڇ���1�8�5�m���%?�:�7���|o�+�ǖ͇ϱ஥��#�"�[���z#R�8������Y�Md��A#g�o���JIH������ʼ���09��ע܊'|�+⥮���#�\��� �2��3�r�\'��q�vK��WÍdfC|&1����ɐ�j�JE g�P�#-����3��0~��M�3t��:���E�p�*�֗����4n��A�o��V��1C.�vI���T��߼��y=���Tx��v?߂b9�iW~��*����l�qi9�,�J�7�*?/TC�j����K�b"��ؿ�عd�7�,��v��!��f�[�* h�{\I�/FlM��V�j�$M�=��K"�;�B���K���=�q���&�SB�A�]�	�-��nu58Y[�t�p2��kZ*�� xj���J�7��.�뻟�8�Zy6���M\z�E��t�9$�[��a�}:I�p�c�6���w��e�\?$�I���z��5���������\��
J�mRu���j8��?��u�M�<������W�g�4~ ݀�D՟��̨�t�<���$�E�!1�q��"�M�ac����|+N��i=P��%m�r��b2���`��;�s�*��9#�:�z]���t��nb/"-f��P`��o�J�}��q�=̃&Y-qٕ�9���7 .����id��$9�������޺�ٚ+ڢ�����L׼j"�0��W'���D�����g)�ڢ���Lo_3�>��#Z�Ր����YM��Ȩ|�D?
���[��(�Z�����������<�%n���rc{�Nz�H]mn9��v[�e��3#��K|�7v�VC�������5�$�S����;��!f ]P9���C��J���6�ڤ����U�;#��*��w��t����u�����J��ݹ}9�|Koğ��DY��N
1�9栕��������/��7��1��@1�d��wD45�1�Kд1.̠���6�D�Ex���j솢��Tc����ʮ��2o"[��4���i�;���G��	GN1C=�GB��o^_d�R�{�颦������z���j~g�[KY4�no3x8>v���k�a��3��Q�'`HR��}�ɩ��<{�IO3��Us��#����z`I�����W)h�%Dp)yΊtJ|-8���O���o�.�j�*�p��(�ゅY�4�%���zF�z���&�Ei��F��=�t���M1!d>&p�C��(�������4�%Ɇ7QDƸG�BjQ�af���^���Ӳ �Y��QcT��Z������q�:5�)�e��9�lQH��Ե� <}��)��@�
���2���V�a�@��V�)���z#��E%_�b�E6�� <������z˻��dA�^�C+�H?s���k�P���-�8��ň���X�� �han�s�p�?d�z>�2���AՆ�j�2��!	���qsZ�Ԏ	8��٪�擰i�.����z�ȟǿ��� !�
�@c�?jh����n�p�D��04<:�+�Q!�j������a�|�ۡ3���Ǝ��C��X��>tH�6��K�&�L�om�hA�z�}/��
,��l���*�+Ĕ����X�·��M5No���P
�7RҐ#jS4A_��?8�Q�!_�s����׆k�\2����|	��5L+�yE����Q���b&�̃z������[9�h���{��~�}�B>�؄ݕ� ��*p�`�B����o���w|����I=���Á���[�c�@���&?�o:e�w�����kJ+ĸ7 i� �����:++؉A�\�wI�[�d�^a���;_c�/��:DC+���:�~�H��BC+uq���*���u�J�[�o��j6�pMǐn�S�I�k�������Y%1��Gt6zM���U�0>���p-R�Dz��b�eI(>��p9b��Q�W��aJquG��I�$�������+l���NF|><o��s}�ާ��T�J�|�i-\6���t=��f�E��V�n�c��u�Z+��7��*�Uħ�<�,1 V�����0��{U����v�F�UC��q}���4��K�s��Z��cI���2�G���B�Ћ)S��@V��q����:��ԁI֖L8�����߸�y:C:�E�ҟL�D�b.�Nc2���/�+R-��e�m;��vW�� �-?�gO/¤ ��;���\��;v�wK�MJ��
f"�g�ۜ�\jL����,��)��ƻ!KP�GĈ�>�rv�J�#:6�7�+V�4}ɦ\����%�އ���;=��7R����#���';,�Ƚ/;n㿅_/�C���M\v��y��Et����?�Q:1�j�3
��)�,a�z�pJ�}�=�'��I�h=�^ #��$P���:��4�uY�$�!b=H$����Di�Τ��_�"@v�n�T��Q�� �hB�>u��Yae,(����3_�����e�f�j�I�r�S.�{�ޮY�]�-�Ye�V�rG�+ɥ��
������)XG]r[L!��9�E��wD�C;*��4�j�a_�ذ2:�(�Z�2g�L��/��0�5������hS8q�C�T%�w��0Ӥœ��@v�5�r\f��jV�k�^SU�����|�Ѭ�u$7=��6z�>>_��^��<�Z	�ze�IgXi�����HX�=�ӕ�_Μ28�Ob7�e�ͫXZ���(���d���{�!��9P�K'�y�R�7�����f�z$���j4,�l%������UC�W1�o0�2��J��s�����؎fM[���D�U����ĸ!�۠Z�'tlO��������}�S�|����*�NQ�� >�x�ޞic�4��l�J��[�)X�w�Ui�8G�˽�BmJt�s�h��%x�HsR�t@v�\�c�w�а��I�5E��i��wo͙e�|�ܙ�8�V?+�(��v^��%�s�G?|D���O��#z��P�����u�ͅ�	�k�(�m&�l���a9�X�Ŗm�uxD��O����!I�|r�^������2n⯥��7r���p�V7,į��O6��G9���`.iŕ�۟3ލ!�j1�Hk�U��#D�vN�L7��%����C9`�y_��Z��&z:����l�m��|� agήKbN�p�&Ev,���Ӡ!�zY�q�F-g�Ή�at��9��3s�+dmC2}��N�:?�N1t�g	osxۺ��V@��I��m4�W3Fl��Ѐ �2�7��Y���_�e��u�=��{�y_,a��csA��M\E%�����o/�z�c�����up�RM�&}(e!�2�k��B7�Q��yQn0:��L��dܛ�^��>!̣�Ӎ����ĳ�QվQ�1W#��qACO������I��E�s�F��)��Nl�
�m�TNs�p�5�"|�'�8�Z�%���K��<>��ѵ�c�i1���1��B���a�;�SO������3�(�����X����
�{�ص@2��m}�/�E�����U�*��/�f񆈊�P���A��릍�ZV_���*��䱞�
-'�GIMؿS�_�}�D����1�W�c�T\�~:��r�/�l��'q��q1*��0U���5"��FU�g���9:�f� �T`|�p���&D=���}�7LVb:J��>r�g�ǣ ���Xcm�o�Q"��H���dу���αI�HDG��zͭ�#!89,(����]����/�.<����'}���������Y��'�:px-�cHC��:\ƺ�/V�.:b(4�0�5ͅ@�eӕ��F�a��Uȱ�E�3�4�jBtא�'����шO%�WQC\<�{�P��[����w�+o#Ů��'�e�agcHegj����=/�}so/�#wf���pr!Hr}H���nI�'BoL�%����S�f�m=��2�2X�:��&0�މ�)���:ᕆ%�NRo�жBZ���b�I�9��53�r;�P�0��4.�G�7Io�#(Yt�P"�� z����Ԣk!�C��Q5��q��
���{Ƀ�n��|x����?�:�@X�ÉY�q��{���ߌlr���|4�?8m�J�� ���I7����ٺ`
��Ɂ���/�1����LJ�E�'=�i�1y�E:����}^����X7�3��5��_�󵯖$$彍��{�T��'2-&_��0�ޢ��!;��'`ˢ5�Ҏ����O������U��U��������c���Ɩ���T9�zM����U�������z~ujsM�f����>����y�&�+00�<�x���5-B|��%@��i,O⑸�?V�vd�e~��9��sչdv�o�l�OYPzP���ъ��熕¸9����1j�b��l|����)��2%ˎ�
���d�PA]�`s�(�	�0`?0sWT�r���"��G;�3��1�g:16�-�S�[>UM�Q������c����]E�3\RmDa��@���3׳�ȑt^�1m� )B�ܨ`��%W�x�@U,���]Zei��dM]�sk$��|���pǘ�(�3ƣO��J���/l��ƭ��� )[o(��lh�!���gCD�<J���b��qtK~��^4��<�me����p6Q��!A�q��9�$�/+�O�"�5Z�0r���n�����;k�g�>�aNKl���ߓ�7�[����y���h� 9�hV�jn�InzGxI�����v��
!'%�h�o��:./��=6|��!~#@p��N����80��RG�n�E������s� �d5?bg��P�k�IDj�tH�F[��e�_�y@�G�jxG5j�]d��%�X�c㈾����n�����lt�Cߦ�	1��M����U���{�`"�������&W���j���믟n7��I� V[$�0:��{sA�a��?�s�a�CM-�;�0Pvo��/voc����%>�)��]���o4��%��;a8E�We��M�K"	��7�G��[���kr#�O"i�ؘW"�ۙ��U��f��#��Zuة�c�p
��Y���U�㝔�GC�8����e/��O��
�c��p���v)@��wG�Χ��tt�/�a��ٖU|R'��
���ԙ0�E�X+�O�ӘB��aY�xq��B������l^R���~ �n�j���o&h��z�p���	Զ0R�a��O�B�t���М�%��.��&[�0����L���2H�j�S.�mropʍ�nr,�]=���u: �_f�e�S���¹�i�XbϛW��(���%�W"���ڭ��il��
����4�n�@-#��ѳ$1Btyv��_s�U"�3WZl�������� �\s���Z[#?�c���%����I�1�Z0��̢��C�,x���M5f��=O�\�Zɑ�����qUn�ޭ���.��![�U<UBY��G�`��+�S ���}}�N5�X!�0(�o��,��t���БS��^摞|��k����u$��\Q�cwZܕ9w䔛i��À���X���b?
�<x��ǋq��A�G��0�>ɒP��d���ŚJ~�?��,(�����\���Jz�v���!�f���<�J��V���2��)Բ�Ze��`���M��?���W*4{��f$r�'�nƮ{�9�����3��5��kP�e���8�҉2�~�B+��Y9�>_�ľ�Ӑ�X����9-���RJ�4j���Ի��j���.N���<tsQ���\Db5}�	�b�4:̃�����@��<�C�]�"�6�{�Ֆ����9��� �j�(VW���)Y�Mp1�����rJA,��J&a3V)ҕt3�{�[�:+��h{��ܝ����|�N]�Ԋ\�E:�dO�-���H�-_A���q!��U�>�����X�Tp,R��in:sa���V�&D�.�-:��ԹF8I����X�1ek�K֣@����wXf���B��O��_�V'%DN �����&nm�,��IjZ�.��Xg|Ɛ�M�Q���WS3��xk����$M<J�Q�
 �	�WO�S�߸��� V�힌�k�6|J�UvC���Ma!45k�=�ƭS���N�j&�A�~x��QV�NCu�BkP�ˑ��D�b׆�o���H.��tETf���o��Z�t�vc�dZg��O�19��n�/�yb�^R��Le�.��#G
� ���B�+X#FÆ��4m���<�ͭ�@���%^f�"D6rz�P��N�gV�l��U�� U�O	��@(�f�@.\!�D-�Co�G���jp~��2p�%n��Yŷ���l��a��G�\�H���q�H�w�N�0��9��\�w�q�"�H�y�Y<����d�۝�f��i�~��+Q�!D��A��	����lV0�� <��[��C6��w�hp�ƞ��ǟ6�`�}jiPq��I�{��.�v:N{I���nf��"�=���j\���Ap��� ���L��lEs�& ��;dlZ�;[�gH�N6 ������nG��u�#{R�04�~���^�J�X�w�^:Xq{�B�Δuu�7J�
����5��-sO��|:�.rm���S?��.�}HR�w`[O�t8��r���=�����e�їx}4gR�&5X�'�� ����Hm�T"a�p��6�^��si�EQc����(L�ō�#`i�A��	�cpz���0�27�� �YC,�劍�t��ȅ� �en�~w
f,��S����)^���?��i�l����t��ݐi��r��9v|�ت�v��Y�,<f��Y>{ؤ[P��A/@��>\�����Ū"q��;����'Y�em�LB�?2����+l���Z�ˇ�B"����aF5��v��6���x�;��n��RE��MiP6�(]}?��D��2~ʶ�M��9*Q�$�a�'�J��C	�m"�v�"<Z�JB�&�>�2*�j����!�A�I$8tAR|�9u�{�@�p@b��F�u !z�8Fǌ�z:N���a+�t̡M��눥�!���	8m���.�sʥ,�Q[N�o�R=qm�5��f27-�<��NC����E��$�0�x|Z;�� ���rg?��U9�7�m_�w�+-*a���'���?g������~�q�s���T�4�+Ƥl�1�SW��E�� �az��o�kLH�Ϭ~-��E/N�k�Z~��|��M[Km��}�P��G���ݗ��YDF��H�l9�צMS��~�у�\�I��|Ǡ�����̎��fy����v��zv�t�P��ʢ �W.M=pڔ��ª��&���O��#�{��"p����!���ws�%�t!��Xݐ��|(j�ݯB��%c�����V��,\��QC��(C[��/����1�s�<�!�h��-_�x^��X�Ų󖑆<��(.�#U����!���S�p�p..�7�=/����r	A��w�8��$(tl�X��10�˭���񚛊��p!�a`�
M�v�`XI빉fr��ڝ���W���q��Tsw��b7,��N���6U�q�tec����G��3)�|�Sx2G���S��U��v���
�qw��*f�3�l�=�HR0��>M���~g�C�d8��l�e߱T�jʢ\�����FR��a�nB����N�o+,�Ai�ܩ��2��pg��\#Iy>r��!��ՄO�_��RK�gQ3��M�sKRکv������#�mb1v��"��@�|�n�m�C)�厱UC�I���������
�2_ͱ�k�G����_d��R���Qi�`�v�<ki/�; S��&�\JO���BO�	��x��!Y_�>�>��}ڲ�I��p:ҍ���!(YS3�s|^�y���Q���C5'�}�_KY���鄯,!J�X��Ѫ�-=%��0�L�X}���ϋ����ؙ2[Y���v��p3R۝�ϵ�#��(껄������nO+�����$�x���e$k��և�r& �*8
8~��Tp�~F����)��s#tб�<_&�0�ZM��JF�և�O�w�"ͳ4�Ha?V�Q��&�3�D�����*���-��;�����&&��}����&ơ��;0��5��˘ QDߞ���+n%���wE!o֜^����f����C��O��?R>�������<��x�8,�}�;�I��e��T<����z�h�+�� ��+)cK��G��Tq�9�b�%g�	~��=�X���P�7�骊.�E���k��[
<Do �[̂i��q��f��A��6G ����	�>�GFhZV����%* �/�:L�5���5��y�)�"�=MŸ:�#}�$5�H��a�[x�����]z@�/g�z�</=�5hT0�N6��.|`�G%R�a\m64L�x�'���]͏	w�f	B�x\����V�m�����(�P�$���$�f�A�4.E.�K��}����� �Q�z�zW�v�h+�dy�V���Ww�p�C���A^I�Uw�%�8�{�&�i}���ow���RPK�W�)��lN��n�҉� q��A��\.o)�(���5�`k�|��5R")RDb�I�1����)v}��<���<��fp@��}Qc��?)fTw����U�]J���B�2Vk�
��LC�	/�1�{��{���_X=���	f�Z�SbR���>�bO���l��,#���q3��J��
�ŷ��0ɇ�#0�$"��~	u�5�ޖ&�O%Ym���C�)M����Ͱ���Q�S)M���t]2��´�f�pu��<��63p�,#q~ʟ���?����:���\�w 'BpCz�,�Rj�p��	ӂ��۳�������ؽ��͔,y?f��뙩�t�e�?�Z�-���s�t�Jֻ�&m�����F� $���,[Ñ�ӺP��,N��J��g�f����ƶ1�1|���3�&3��ZO�Ɔ���Q6|���gq��I�+]�e~yr�c`���@rF�j'H�!zr�4��<d;Z�Q��ԣ]gT_%�=�VJ'�AS�a�Yw�XRo���6�>��6M:I�:�)R�S���*:���W���"	m�E����TK!]�J�ћ:�����"Kv���m�OC��O����1d���S�y��-�*�W�E�T�y�b��mB�j�������͸�Y��MfݩCb�Rg�l�X;�rv�Bތy��,�0��#OI����>u�U�|���0�(�=6w�u��	<���
�i�8���gp��ho�Y���v�zd���P=A
�ʀrO�f�fǐ ����<�x��\
��\a�l������nN<%��uź%/Y���:��Ry��Ӌ&��0ۥ�B'F	�56����!�h��V1��~�Ϸ :CT���:3���>}Xt�C�Ҙ�]�/���9FX���$n�E��ry,��;H;TǾ��s�A�6e�.Ma?�9,�]�RM �	;i�HVD_����h���ϡv�h�+�����M����@V�"\s��[l�5�����P�p,km���)���X�ȨF&�AK��t]�Hc.��H"k?�����K��M�أ�5ˏ);*����쐰�R)�MN��2N��z��~��H�o�*y��{3}ms-���toæ+���iF~�h�j��
8��2��c ���q���2���k�"���6A3ΌE6Au�ٛ�mk)K�E}~����5��U��9vsN=r�Iz���o�{�A:ezv��������=��	���,$�H[a�1b/.��t]��o!uFH�4���)���/W!��EƘ��Xs����£�N��OA�?^�8+E^��Xf��}��Imvn|nY�`bʹ�'#"�ӝ-���u�L݂��у�G��;r�F�E���`NS�P�s�-Ъ��&o������O�m���m"�_>��ܑrc�6 )�-�-��:0�==Е�◾�����"���LQ�@����섌�:la��/!N�㺪��k#��q���P�$�T�&�+�5��z��Z��C�Ye�%9��R"�В�A�I��̶/����`k0�
"�3��㵫�P��$��U�1���p,�X�G�d�3˰q���@��e#$�Uj,f��6l����.���'�U�=?%x ��ܐ��;0xi�O�B����Ҫ��Aj�u'�R�� 	���*����I�C;	L�A���u��|!�@Y��cj�c�X�>N�o�",���U$�ƮR>e��S���Ψ�/uĒL�<qP�����
A���C97�D@�0H�^9��up|_�7��@��+S;S}�^��d��w�Ԋ�I�/Pt���T�v�Y���!�E��Oo��X���~&DwOwDc<��CU���?4�=�H:�5|tO�ٓ�0�xÿNjd�/�s���ʿ�d�~6���)�	P��bo�d��� R凫ڿ��1����uX�3|�0k㪥��x}.N6@4�\`��`������(����]Ӣ�ɧ�$���Z݀�K_0?EB\a6����zzn��_�����{��	����5d���ԉ��:�q�h��t�q�Ҩ��f�p�G�6���$�y��2��4�5D[�w���B_/��\
��^Qd�kAy��6D��c�p�酎���
�a�)/�ݪS�s"��Pj}��ַ���Fc��U��жW�l��[N�6om�ї�wAF�ńE�L�9�����!�k��i�E��겋�ǘO�iK�s=Ѡ
r4�{�/d ����"�[sK�
!��`p�RiY�����M���E��qHnjS�91�jB�^�@�:�O�RN�[�>#��S8��.>"O�~d��$��0��V1^JN��6�o��ur&�"���+ф$�����:pA
��?\���*��M�M�O1J��)���b��şm��1rPxᩬj(�
ݭ�ý����etw ����pXq0�~��C���Hh_�E��� ���7�|��
�Q4u����j/;�T�;�s�6!+���WAk�3-Z"��ݻ��\0_�Vk _���~��9�_��Tx�m��k�*\�6SP�_S��!I)�m�*ɃG�Z�ݒ�����|A�	��YP�[c>����u��	�Zg�`o��E4Et����v�a�T��𻅏c�4��P#C��$Xw蹣m��;�[����[e*���vri	�VKE����Z����JVU�On)��;���z<L�v\7�U ��.i��?�ϗ�Jźz���:n&���6��������}%՝�����{�ˬ�vG�N�,�ACthOC�{R�7�CmN��9�(VS\=�����`.,�F��Q������68R�%�V1<^v�������V��V�M�Sx��a�`.�I���_�E#�	��"Ņ�.��lT��Tٱ� 0��5ɱk�~�\VV�0�Ɗ�����
kٟ�m.ب�v<&%�(3�����D�l�k0���5Һ�K�Hь�d��
vBT�X4��zO)��9$vK�
�U�w�O�5�(@�faP�@�.P��>(��f�G���0�� ] Ă�K��-��tA���n�$fV�ɱ�a��|�KQ�!&�_�*��,l�����n����Z�^ݎ����� ��
wt��L��y�/T~O�:$�S�X�wps|�>�a�-k���94ۡ��bs�� ���I����0n&ɉ��/=�X�<yL�X_��JBat�rj���&/t@]�xw������XEXi�Wx�llJD].�s#�;�~8?�vXG�7���[pk�gҫA�ia�+��Rq���t�g �̑�{�2F�t�^Mj���,�#��Ζ'<�bf��>'�qFw/�kJZ�����3�k ��?�����:�(@��ǥjxY�M�^�}�=�b"���{zeh���cWAP�2|�HL��(N����e�aq�\�g����d�V����i�v��gͫ7����J#1� a"��ځ����	�I;n�p���A��!���D��knT���ui�r���5�Z�����?:��G�tv�,��h��Ʊʡ����B� ��D5n8eJ�[���v��O�D0���:��ɧ���.烏h���V�P#et��X��<�AHu~�1r��[0R��S��)�]�%�-�!:UVm���>P��U�����Y�C����R�R\�l���=U׼��KTr��	sf�L(Ơ�����T>پX�;�)�:�yhY�Nɬ'�2ZUT��A���ԆIɍ��B���&)�i�
#{�r5<\��ZQ(�,)��чK�� |����t�tpԺ>x�N�0�&?�e�R�z����=�4�N�5��}d��k�8��|;6$�3�I�#yؾ ��H�j�%����É�xw��P>�G�譵�Dy�á0�����ˇ��$��.�(������]�[@�*����{��+�eh�C�S��w�f�c�3������/����8����� 0l�"���O%�%�pO1m�#<}�
z�o��b�	uˉj�Z@�w�j�HV���TwR��ZC���c��{�㊱\�̠({�7�V�5���7O���Ӂ�ع�t�xw��M�f'J�p��	������?��������ӻ� ;�AMR���z>krE.��E���_.�C0�Bw�tl���������[D�^��O6䉿7�-�ND�`���Ht�V60�b�s0��dѴW��W����`l��W+n�q��J��PT��������������*D@��ʅ]���,j&n�� �� *��J7�g@2� U�$w!�qHM����'��{L�$c�����Ѕ��ؽ�o\�M�4��4g~�'SL��A8Q�ai' A�I����57s�x�69�*h2[�U-m4z<������J�"�ؠ9���1Mod���&�����{�ܩ<��S,��:=��$�3���S��aB{��ʩS4���:� �8i��Q��8}�;lK�l_��y[W!����� ;�hK��V�o+���I C�D����c(��-�H������p���������a�;c�Ϭ#nR����W�j�CIL�X�xEq>'�q֛N>�ă8�Ӎ��5=@�E�"�qG��@��.x�dU�1AN�\%�%S����u0c�oSC�u�km��u���8��t�Q��j۶g�cM�C���q'���}�ē��uPX���G($-?�}�UI�t��1��w"j�1�t��}֮���}6� �@���k��![�	uGN���zT�L�O�~1i������1��2��(7ya6�p����v������|�E�����t���ay�vlS����=�>¢�t�MF�R�[��х!"�NL�=b�n"RoiN�+�|.��e���������# '�w�"I�|:�?z����=5�[ͻ�o&�r6,��-C�7�2��I^����	�f�L�7��2��i/F������'Ÿ��~	�
�Z��o���r����M帟0:�L���FG��J ��������������.T{�7I�t��Dq�ǅնM�D�5�V��2�x��2�g�m5,H8�^�7��Tm�]!��.w�2_U���g�R�	��΁^� H���K8�>%�0/�����u��#��&+:��A���`����aCÉ��ߕ���5]�������y�@P �x2���B��me�Ӂ�q
)�~ӳ�ҫ�ױ �4g`�� y���IRn�꘹���	O���p���:��T'/-��Leg;���R4�n��X�UB��"^�
2v?�ldؠ��9	թT\ti���7ޠ��6� XSP�e0C�!����uOn���{�Dkq|z#�Q/zL�Uᖅ ��WHK�XwY���58�Op8��P��FOx����^��������(2�
�h=��"�\T��r��
M)�[����:C ���,��$��&O�E�!�R���:l�O=R ���S"� :��qҞ�9U����_^zY��������G9��?J�Oj��^��,�Q���b�6�XJn��I�mZݩYߡ���Ż�{�a&�+BALx�����~������8ʥh��� C���8��2��SMrO>����@L{i�E���4N#R� 3�RѮ����`�h�.��F�nIm2��,6�eu��d����d���O$|��#��e�<� ��4�&�9�ܶIL(���۩I����G���y��r�lBl�Ig��]����3��eQ-�N�zg�p$'�H�W�h�b��~�y�ױ&`zϐ�dx�~8]���R'�܆��Lr{�}�e� ���ސG���4*:m꛴�7xA�So0N�Ls���A �W�8�*���`wx��{���C�#��l:<3t�Q��@�|�q���'�A@���<S�Jn��]�x�ӛ���H[|�����-	�(t�ҋ�CVd8�����҉�ا�����v�*��sY�M�\l(.^�L����i;�3v��fI�գִ3[Up�������^�`7'�"͌3��C�v�"rj P�(��< )�l����7c�a����)`g�h�ዴg�s�wڴͨR��3��"�!�ؘ@��~H���o��S5�U�7T�iM��y�wGU��<>���d���|XbftZJ��� )��>m���v02$��4�^�J�\Sa[vd,�y��.;]�
����Z"�j�{����(��Q��
�����S�cvx�Z��z��iHˠih5e�{�����m��Sv��n���*$�lo�����=���G��|�����Ve{}�*⢱��~q�bx�4����E�yv����X�%�/�i�,б5Y@I��G&}!̻bL��`�oT���~$t�5t��t��D<�̱�T���w^j#@��*��R�A�J+`�R��?Y�E����8�TJ�u_Of�����q���U�T�c��M��6ߍ��BL	%�޺^���S{Μi�q�lW�x��x�; n�g�AE��X0����l�iVTŎ>?Z��y����p��Dk�óO���Z^Z�	o�_�eT>�&�f?��' ��2��*&�Ul��o��K����(�(�}�s^h�"�*l���L-g��&[/w=��'>`ʐ�@�UM���0+��0�d�*��7��-	W��e�T|]�,n�-N�5Nm�����a�1AC)�'/;���#1�`�T��2�$�Jqb��D��n`[�2��D_��)j�vӪ����C(i� f���f���
�V����X��0r�V\*�1�m_`bҥ-�,�)�չ��ܐ
!��/�D����@:f�c�&-��:�������4>�L
���0��	Ȓ��׌��20�����) ji�����s˨#��z�"堨b��%��>��x%���y��r_E�t��SmB���k�ۋ�Rw(M���w��y�Q�\.��y�4öZHnB��EY�������ԝ����&�����)R���6����C0	I��6ҘI*�`�O����Y�[$�I`�!Ÿ�E��3��bZdQ ��-e�C;�ʊ��� ����b�ޔB�0�H�vY+妲*M���,^+2�����0�jI��zL�Q?�=�o©_��y�M�K�[��4�5+�Hq!\���q�������q�.Dw���AAS�;��30�wL�c�̰O�E�8���n���*�\�'�L��C��Xγ$�w�<�(��S\r"�Q��j�V����!t\�"��%��A55��)7^Hgc����s�M��k��CF²Ouv��i�&�o��\�#˔j�_�/%��]c�D�ۼ.���F8����Z���~A����흰<���<�}���|[�Ʀ)���;$�e�U�r@�5����3�|�������w6�ּQ"�9Kʤ4J�� ���I����I{]=d�*���v�V!���L��E���J�X�����.�D�w�
���׵?yH�i���~�R|}=p����������Q�_�?��u$|����F��]���
q潐o��S��0���]1��\��Ag�7T���q���LI.�)~�㧠3�'ͤ �)Ju��v�|��7�^k�I,�	�o�� |_cwW�
���*�P� ��@���j�w�|��@���D�C�v��s�F���\�1K`�_ׯplT���tMN��q����'�����z.��/�wZG��r�ٜOE��5t��=D�7��1�{���_G�@f�XC��S��9��ցy��:Iy�0Q���z��]c�A���dB8��D���TƼ�;�Y2X(f�4����]����0�f���;�Ը��rm�?��:�Ӳ�B�`��(�'�E��P���Z��扽P���]N�$鹠fH��^W�S�9$�u� |���[��zzh6��K�!,�A��c�UD��(����^���q[��'
����^@���˱Gz���{��[>�R���7yЀ��@G᥄@9/s�Fj/�+X�+j_ �sf��7p���X2����W�� :V:�
[d��ׄ�ϫ�8�����5��|lY�>d�2ڢ�+"7p�G4.���yx���4Ó��,���U��5�a�6,���}Rm��c!"2Ң�冧>�UL	FSKF����\5��_���*�@����.���jZ̒3�e�=�_�0��>r$�;Qy3Y?���/\�qH	\xrs�	� �ܭ�[e��]"�*�p�Յ!�,OzaY�l��D�n���$��by�/�5u��ց�@�
�W��W$�g+�Q0�[<��e�������,��4�wW����ks�����K<=j�@��ƙ_��GKWT�td�x-�:򄺏����O�z�ģ�.<����!J�9�EY��'�5�MC�w�!��[�p�6V�e�%�j�B\HK	�x^Ӗ��w��{��#ϡ��6|�:C��4.̿<X'��S����8_4�3�c4�Ҡ� } YTi��!X6����(�����KU�i���F�	�X�|3Wr�͗�U�����L����"�%_=���G=8a�)�b&�aP���-�JIՐT���1��J������,S�9��2��n�a"�5\��&��jz��^���j�G7���z��n��u��l2K����>�3O��� "��`�w�<[�23a@�i<S�j�S�ES8ն�s~[qa_ĺ�/ԑ�k��l(D�˒�т�$O��iY��m<3����=�ay/�)~u�ڏ��3l�"/��vH��I��ۍ�r����ڈ�Ke�F�`(��LӼ�H�"juiA(٣ʜ�Ib!����"V9�}��Ҷh6�7z�t�Y|�R����h���A����]	����)�3t����?7U��|�gV���aA2p�0=� ��`��%-{Jʜ�:�<do��*�Ņ\(��#}m�T( �\Z3���jp��I���AW<O�x�nnH����
C?>#I�Ey�����(�L
ѷ�&��8;�9}vW/0�}+ �7�ZRMo�9��=[����#�;F���<x6��f����Q��`ڊ�S�i���},���&����Z����jB���(�8�V�����EÇ�\��TNn�Ȼ)Lx�K�?�ԉ���X��z�xS "*e�g�!lw@Fu��xܩC����ne#Ya�Y��DF��� ��=s&��(�����XUk�,�V|�r|ӎ�6���!z���D-�	S���#,�S���6�F�Z8}&fmD>>!aҵ0�(��cAu��wI�c.}��p5b�"�"�b$;FY_E�|������_�P�EC}�Acs�W̎��8��.
k�"|��l��	1ֈ)ū�^~��ӭz��n���MYx����2�<�V-���_H�+�4p!��V׸^���o��^��Yޭ��.��NX��म�m�ÄD�� ˅�<�:=w�7�m�� ��@���F��R�VTru���;���>+��X��q�,,���NC�]��3�3v��B
x�n��E�Ս�|��	�l{%-ׄ��7u{e4�8O~N����Ku�4�Y]4���@0q��AȌǍڗ��i"��yjY#����(".K��Ύ G<�"��ހ�����@�����9���%�2�V>,�F��T�.#����6%v��u�������qFaa��8���5��'�]�7����4��2sy`�KZnɔ�z����L);,�tt�X�Bj�� ; ��G�5��}��d:�{i_��'�c��+&ۉO�J��
~�6���V�J��?��rx��j��%���)c�t�~� ��ڢ�D�O	䧇�BRV@�����8�s��U����}��!���]�wfèv�yI��f�O�,%��vQ�Yv)|�A������n��1�q������ѠJQ]a�[-�SZ�=�5Ks�8|�^C�/��;���ߊ�G������n14�t'��U&���C���ZA�<����%����ÿ��LN5��N��&.M�p����;{-�i~�Jh�l�ɾIt��p�_��ph���5L�3:t,�L��E˘�1�T�8ͮ�"�MP(23��,�? &�JEk��tj��]<�~�;E���S��a�PkfJ�%6 �o�[�n�Y�I��B�fVj�Z׎N���^�w������OG%%�G����f��`���$�(�0<g�td�%`9�n�O��;��̄�xR:����C��7}���S|_|����`�"�����í�^ɍ��%逮PV�jR	Y{^B���χ�j�+��=@�)"�Gx������E� g���_x2*e��@��E�2b��#�w�$�zW�j�������E��N�X�c6�,�b�`�|����	$��/�YN�����-�c����^֑���9b��o�i,Z:�kD��&�B,t�R�cC�l��i"��rig�����ޠQ�+�w���յ��}��L�/R��aNj�2�_��/��1���%?�SNQd0��ɓ�wֆ@��C�=>Cu��ŻKV�嶹:�:�i�tH%������+ӟt��8�
����-$Ϲ/9$֕Q�լ�Q�P+��k�����﹂?�3�7�ѝV�a�ҘS����ҵ����� @eL�>�4��B\�����)��t'��T�];
���m6���R���gU���|Tuh;����J�dj�ǐ����E6@4�^v�D����U/@��/���DJJ�M:�4 ����Ԟ��Y�g� Q�5a�k��x���"3.M�4n�e��Gv�\^:�i��n�]�Sw�[	x�/���k`� �ek���bB�YZ-���v,�u�r:i�&��jxZ��~��e�sN��E����p��p?q���`:�m	���El7nCϞ����Հ�fF�����v��g#wdpr+u+��r�ݦ��2#$v�7+=&Ap����X@�ڗ���9�."�>)M��-��?E��o�j����ҙ��+�,��^ٮ\�w���̯��h��3�b�@�U�|'��F[�|��u,��c���-��T��������w<M�gL
�?�Dc�˽�e�e���J�/�T�Y_I��z���&ߟ͍?�͚Y��Q��wL�~$���p� 7Ʌ�I_$��<k1t��Vt�<�b2��}��/@29	B�ta�'|�0�q�!��r[�H�0����I�jd��i�=G&}p�'��q(s�*�>�G��ΨD���z2!	��#(S������=<^�|U;5O���L�A#�H��Ko��:�-�a ���E�ky;��f�$|�h��[�w����[�!N}G���B�R��`��[�R�I���?��!�26*�v]�p�#$ ƽ'i���U�vr�{������n1=ږ�l��Q���*�i��s����({��x�dvPC�a���*L���TS�1���>Qv����f�VM�f�5$s�
ml�-��q�F4j�GG �5��E�����(�VF�q���5��HJ��f��Ï���2t��N�^�}�ޥ�X ���>�{r�O�tU97*h��X牎U(|&��n�[o�i>4\�������r�	rj"�-���2{���'=�����Z	�:|��<[9n<Ó/��;�j@�Wb��V�<+������7<�(x>��/���8!Jw�2i� :`�B�I6�
��T��F�T������#l0��5+�ܮ�\��at� ͇a�ƕ�*�
&�3����Pf �V#� ��Py�x6>�^8홮���W0Hه�UpZ4��n�~3Q¦�r��M�H�|���_�+��+��1�ҋ���dI����D`�|z�xx*���s�`�{����H�9�:m��E�jȇ!χ�΀�|�C��)��`���>��)o����2��� *��Ho���Ĺ�1�U����9Dv���s���,�KG�k��-�$I�d^��1�S�F� ��ۍ��Ʒɠ���4�E_0a��p������}z*mz%��\Օ��;��g�>��MB��K�J�E�n��!#�c�H���2'Wv�vK�~������"��L��W����C�TN;j6� ���d{��j��m)�Q�M�>������5�p���6q>b���s�=�ӥ��a��P��&t��nf-����h�&iq�Rߑ8̸7<Ð7�G�*������B�O�8��~0)zQ:)�H	pٌ�WEBY�`��L�m�xs�Ԙ@��"�PXg\�W ՝#ic��8%C��
��$���Ӈ�zY��xo�kP��v*l�4�n���,�6<^-!����Q��@�e-������;�'��s�m�X���A��%�"���Ͽ����r��P)��kg�P�-<�Jv:��h��w�"��`b������[p?�o
7}�g��_:�[I�b<�SG���%�����i�ދ��-���|��<���0%Q�T����L�K���	5t�,M�!g>̃}�n�Z�ՍV� ��ו�+�7���<�	�l��R���m���l氳�-Mf(~�C��pܕ�(Уv�#��l��� 36��#�y�t_?u�kA=�Lhx�ڧ��N����d�����Bէ��� ��ý�D�=mm~�ޥ|����F͆4��H)3�*�9�6}_��;�::�(!
���P�ʟ�rd p}��0V4fi��5E}1��$ϱ�/�&2i^z�ڜǂ��t�6�v�u='��uw����X�����A��"MIQ9��9L~��X��tq�b��42����֥�=��QJ���	5M����!��Po���!�}�,��� G�����\!������h����;4�b��F��hI�c3���=��Z��B�j�vR��t�I$����H�R����o�r��wd�=�
�O9��nu��7>�|O�@�Y��cV�9h��{ �]L�IcR0{��b�*v���)��a+Z7��7Fh�k�E-�=���/�f�*�4�6��	د3��֤!��+�,;�9OK��U�1�.�zT�� ���{	Rì�5b3����:����(,���B�-_ȁ�e�5quv��[(�Q�/+�;��V
	�mw)�+��ne�9�s3�D�=�����!��'���#���W�)F[-Z��?y��kl��D���/(����H���� /���	�G���s@Jߤ�5�u�d�_L�Y=��[&M�˖�)�@ߐeT�/Lr k�i'�ߟ��M�oTa��;-��P�i��Ar�����H�eľԽ�.{2����il:nG��B=�q�*�a�ϕ������>6>ʹ�ۓF�f!�h��Hf��z����/n�'36F������=�8�蛟чjU�?z�c����L~�H�O���Y�5���B����4�6�	��<�U�!�m"sC7���rp�<���P����b�z�1�`��<�o�/�m'�N��~��p��n	��!G�ΙRA�B� �)ە��K<�5s���w��{��|���t�+��a�����i�i��-�cD��<U���j�FkR����0��@X�Յ�^6*S��/b��Yd�g]�8�/A�H,Tw�0V񯎝[Th���4ѳ���hqAs!>!��v6�=_;��	�zV�a�a�/U� ���YtX �6yY7#��p{w�V��B4K�9υ���P�KUMc������:��H��{L�(��iuqC��Դ�nŽөT��q��'�|~|��7���I�� m��x�։�&����&a��0����SM��X�/L
��:��O�q���lȸc���DԻʝ�(��(�L�du,W_Zx�`�\;�;�5 ѭ݌$ ��]��*�xT� 	��޾�7��oSE_��}B�>�8�~�Eg+P�$Y�J_P.8�K���\���/ll��ד�p9D3l4(�T�[^�U�H�T�H�+��g��V�D-a��T̈�4w6bA�R�-�X�����_%����]���h�D

��v����}y {�D��a�̪��dn'�4d?��T��.��O�Z��$Ӡ �l�C�e�>ڱN���]=�nM�e�R�˾�����hoK/3+�g�(5�[��=L~i�(|6&Dl�?��]n���|x�ñr���2��p�K|�P�y�³����}O��f��8D��SM�+�Y�4r_�c*� 3�n�l�M*�0��S!���tj��I 6T��AӋo��.�p��0�iX���R}�B��Qd
�Zda��˩��z��E�r��H->7�G���bV����K���u���� �Nk�"�ʕ�i���.�80/FD���_���<f����S�8<�Fxyy�ٟ>�Ŷ�
���0�e�'�����u�?À���݆�{*���Ŭ4Ȉ9��u	���ʠ�����]:�w���
cY��M�S�����\c=QEN:#�Zn�����;���Q�5[̔�Q�Z]w���D��}^�ǝp��&�XNʎv�)H�6�	��8��Q�F\n$�?+��C���%v�^���듺�e���&�� ��*w�T�
�	6�I�����f��O .E}�z>�Wk淁,[]���AT�0�&��°�36�T��&Eп����F��4���n.+k_N/XE�/>�A��ө#��w)0t֦y�6����7�N�]A�_,���<2�r����X��9FZ�Z�K�Y}��Z�5IA]�/f+�]w)�~ܦ-�H�#�v����x23�1-� ���@��	�ӳ��6u!χ>�*�;M����{�;���+�8�@MTzѹɟ����ɀd* �;�Fv����x�[J/+�kRg�����X��怒����С0{%�z��(��;�_ç�I�\ShC�h�&�Y&��x�h���Ϭ8�.��{p�ZOz��&Ɉ�XӁZ6ڍ
@Uh �Ao���rC��� h$W��t/��3�O�a*h�jU9x[JI�P���{t=�yYm�	̩���уp�q@+�\M'l+���>�ˣl���R��ͿX����W�.�ș3g�Z�7��� ����\�u�(�W�*�B����,�]�j�t' �8��1�Z��I��Z��̚$u�)K����% Yy�t�мM�<����:�~CM������麭A�����G����δ�je"��0�fDs9�R�,v��]�x��>X5�\O���I�10[4 H��.^��g���:SlI�f%(�����!O��u}��g:��د���,ORD� �J!�}�#���LZ���nNOZ���_I�Hiͨ��o����}��q[����%������˒�����*���&N8�A�0+@c�Řp������a���5�Y�`{�vOb`	�icG}CW1�:��
����)��/�k� Tka�fFz4�#�Y� ��n�����l_��}�O@(��;���s�qx����HV�Hj�𡄘[^n�ZG3`	�rƪ�E|$�p�Y	����cl�Z@�L`j��Z�tk:�����r��$�}�A��͗g-��@�qܒ��_��-,����'�ɋ��B��*�'r5��ِA+�P������TuI��}�^��g��he	r��D�=Ua@:�_v��}���<�b�U+;��U����_6�N���«)7pu�[��EQ��]�׆�٦3 ^�����pYV��xҌ<�p���-��Z`|XvG45ɤ����bc�l�>g�� s�7_��%�R\9��x�����&j�}9d����Q!��B#�Aj!�f�y�ϥX[;}\ϲ���|���j�+�T�p���b���E�}Ļ�h��
�ȶH�4~ŊZ��	���R�{*������D�2qf%�wF�i�A�2��ٟ�rhv2S���d�]XK�4�����-�Q��)bw�y�3�gz~�P���nA]&�@[�rZ����6�>�V٫#��e	b��� �i8V�_6PԞ��_����X�ŭ�H:s?
7��Y@�sA(�	��
g���?�H��"���Y�r�᫄�����^ƺ�s(���m0M�I��{�d���v�$?{O��[<|v7�Y�/~ɇ)�G�J�D*���;r~q����rة���c���FNf�aӺ���������J�|uX��]���Y���5�̒���Uf��"Kֺ��ײ���F�z�,��4'e�|��d�x �=����Q�{�ztb׶����ʳ����1'eT/.���ٌy�0���_LFݟVBY�_v�"�a�2��&Yi���/¿����+:驝�x����c̣�CIvk�47��>�1�l8����,�*�O���L���{ֹN�lÄ�d%F� ¯+���'�u�Y�q���/�0HtK;�S��O�˚u;Q�aϥ��.iU�-��Z�x���:$�GOMj��FK/~��=��v>�nb��<��k*��+��8�8��+Dt��5�+���Ω|��T��ׂ0g�g;�l3.9 ��s�?*�#��;F� ������ ��@�)�V�D� ��#��p�
IM�����XX�1ﴚ+�X�bp_S�Z���N�%S�4�n�}�:@aburO��%�r��ڧ㯩�Vn����,\�h�1����r����Y�!n�z0�_	轨��g KZ��@i�α�%��#lX A�L����T�)�D ȏ ������ ���'��0+����Bb���K�7���%o�U�bw���ʛ%^��{�W)�,�#��ޑ6:(r�T�����Ӏ:#c�رVR����:al[�[C?ΐ6���4�'>������w�B�V��X�Ӽ�<����0���^ᕪ�\E�F>�rWy^b\�U�����j�p��$��E/� 	c��q#�vԺ�`yڧ��6H_V���`_X�z<q��(/B��FY$*F�	�z�0�kM�9���mcP���$��p��TJnjt���s7Ǯ9�3�b)�V�M
��������uB₀��)�b^�a#ܻ�F?,+!j�H<������*���$���i��W�zT��w�����PFk��E�v��Mtv��[y�����NNX}�jJH�I��.zj����d���푙�s{���]�� ��Tf�v���6�v�y�@�H�y�zu�:|fKh�o��W���H��E��<�dS��ϗ�a� K&��Kr�E�_L][I�dA�;�/*����;�&Z�,�ni�s������/%g�Q~#��;�8�ԩ�ǣ 	ks����N���j=O���L��+O��L߮YF'όM`��'26��%��K$RD�e�w��ܵ��B	���ڴ� 荒�h�ùmF�<�(N�37���Մod�9���-��T������@׭ⱌ�UA�T��̮V�a8\�AI~V��D�{A��^��;VI�1�z%��c�6�F�
CP�v��H>��X�~/����*�6����eo���K���������p�"^����h.)��/��\��M)_�}��X��W֩-mӈ�2�s�p��X-�v*��ߧ2�~Q����C���K��.ֱ-��-KQ1�7��^����V�'�>?�9��h�Ȼ[N!�uǾ�0�k���n��3	�B���C`/�)�:�x`f&{��8¯��_;!��R`��[��w����E���-1i�h�I�x �K0l���5Ox9��'�K�.��rW��L5TZ1�ņ�ivQP�"��������G���Cc�R�UY�<DǄ �k�]�Ho2�w@o�IC��1�H_@�VI��+5�^�Lĕ#=
`Y<��p����[T��_������]��'!�a42sO�Zcv�C��kX�"v��^��<gF&���k'y��o���%�OP�Sw ��fIevg���Y@�����ZA<���̱Z����E�ϜO��^fY�쎍�!z�;C?p3����s���s�8�S���
��Aa���Z�W
�����e��U�>~�he��A�o�5]�L�4����	D���^`���I%�L�y���J7��W�3[=���k�RkX�Pj��c�+��R�!p A�*�VfLQW�FH��T��xFOԇٴ�Jf|��C�@yd��kݎ�ƈZZA�x����+R��Z� �8hG�9��%��CE�N���k�H�X=��̒��qhy�r��C�� �:z��#D/9��ζ��
b}�cr�p`>�G��=\�S��R��]1�"K�4���\�_��	"��{\�#��i��8�K���늕�Ws��B���>�{���	��(�W�!���S��TVv�H�o���n�\Um�1����	�{�v��K�.�=��i�����[):�v�r�5aQ(w��`��U���%Y���mng�c�kG���4�k�ľ��0\	GbR>bEj\v+��\M]�e��	�(�Z�1����D���F����zOPe"�=������R
��w�����5�4��e���~���1�x@n�r��R��-�b.y94'I�o�2�O�pR�fyH-���7�M��7	�����3�Z��k~UR�{�i���z�Ey�z���jWF�[�Q�}MI��n�H��<�z!9�0�.�Yi���@P]���KTIii�c���ɾ���,��A�p���qm�O�~�MG�k��g,�.h| KǴ��Y3�z�%K��ha ��aQ��C�n�N��F���\&^�3�P�f˾ MŜ~��	�cG���O����*f]�q̦O	O�ۨ�D�T� �bbF��ٰ���v��KiǛ�(SK�rS�,�E�4�U��R��ƪHt��ZFop�6h9�﵈�
W@d��mC���EQ�		.��D$�O@�er�����{����hM��� q����=>,/G�ĭp��\�)�4h\��G��$�#Gdob���8PL���ZS�K���m��F%�l�І��R��C2?ԉ��]΃5q�p�H��sa�o�E}I�9�2���� �"{QU�y?��X6^��BD�nLy;����R؃���
�Zf�N~n�|�I���pX@��C(|���%w�\��z��O�YOx�f��ks;ŏ"xe�͖��y��`�b������e�
3;.'����\O��ֺ����R����[��Cz��Y��y���<x t#�hw�H���9^�LS�v�,���.�����N�=[��3�V��o�� aa~��ITS�A��J*O���Z.y��!Z����,!̇�,Α ��pKJ���N;�hQ�0�n�!���fp����B��N������V�|���s�{+W�ŵ�Q,*��#�(v���q����_o��	hޓMd�e&�Gu������x{�)��c���<�O���
#��5;�mV�0T�x�����9	�sU&٨������/i>�E�d����>�ɐ0��c�j{VkK\Jz��~>|��|5S��/|�?'pU�ǯ<`�1<��A�4���� ��Qw���4�g�?u�X��?s��G��_�）@\������q	!&��P)!�m8�]���8Hg<*�D;��;�	�0�� ��J}8-��-m�ٺ�,�D�r.��,�������Ԏ9|�g)��Ԥ��`�Hk�S_.$�Q��0D���V�}�������0���.ʷ��	*��-f?OR�=�ug@���$Б��ʭ�B=BM^�wwxVZޫ�,u��J���*A�ǜݰ���h�<�w����fZ��>m_!2�"�����^ͱg1=:�^zX�V%�����;v��{`��Tu-B�����C�ĩ�m������}ǘ�$4g�]���� AQz�.X�� <F�=�%Ә|/�mE� !���7?��f"/+D�#ZQ�v�:<�����y.ȿ�JxH�U~n⸼ 2����;O��Hh��C�h [9�,G�2�޲{�+�ts�-�9�	I�q�Pd Ƽ��B��p��Y,���?��yv$�����R�O�����^�?w�#�o?ܰ�A~M�>�T���<uO�:��I�3��혖�X�3�2|��#�E<0}�����,)�y�"W ���ыm�H3�b�>�	�)&�Z��_�>��T���c��J8p���0)@��-)&:�i5��z�YA���1�^e�/��}m�0���3���ٖ�Qn(��N����ߍ*�X�@�s��W�����g2_�I��j/u���i�S�'H���^�cɻԴ>�#���:�1�����- �^��}���2�XG�iKZzY�\����Bhjzn��=9��TzZp�v;�S������B���������Q[򘠸k�5&�����z���DJh�F�l�Q��t0���0�U���ݼR3���j|��+x�|�@�����|L�La����	��� ���Ŭ=P���+|l2���H;���t��DcjS��Ʈ��	 q����׌�t���3$i�"�voV|�tR{��\�^�խ��q��*e�#��0@��xTǋa�F.>9��딯�;$��@�ި_�Q��%�#ܚ�ɞbu\x����І��7����9/��bV�yT�ҍ�%�[ �k�@�Q�m��D	5Q���DcN��i���cG�\�����3���L�4�����^�C=�tgh��εg@���g�Q=�!\�C��:�\�߼QDBu�[�~|R�`K������I;��|�U1���\���HW�(x['���\&h���);8�@����|�vo�pK] ���,�.xR�LZ�r�Z�
ڔ�Uu�p���/b�[�]F�	���"�wfSIkB�,�" �*Na3]�q��,���G��nb5f�L�B~("\����| J��YRN\�*�����{φ�n��qR�E�}MGj�1u��Ω��*�
"��:�B.���( P�X���=�k�����?khE�gUxp����P����`��q�t�'9��[���5u��U#]Qܵ6�Ky
����[sJ~_�u3s#�%y�����֭���I�X�,���G��ܑa@�="��%t�P�垈��s�����v��_eā��NzJ��3��ֱ��@n�Ñ��oLA�,��G~���5�>i)��W*`�a3G�vԹ��ξ�e���%\��EK~4��ֶk�u	%�71��a�M�NV���Ύ���U��ܒE{v�bGZɋ�������������W��7��% �����e�N�z�����I ��k⋫���w�g��<��FC���v��_�I����&b�pg+B���yٳo偂�X�,�PZ��k�8����� ;�g��oq���+�ی�Ʌ��\I�tYs�V�ZXCT���A��_x4�=��8ҏ�j��F���ω�ۅF�W�����Nb��=d#x8ݾkP��!ԏ'1�Wт§.�/%]���ɕm:��kN(�{K<���!v�
i0�!��5��ܘ��"4�G�#��s��r7��]O{0��[	����V���.�z'2({�/hZ��LF����n
>��{F'{��_N�����g��$ƀ��X���a��]�)��c�]�����'�/��l�C��~;.a�Fm�3����:[�X�@/�x0n���9�\8%�ع]�f#�ͦ��yv�d�LE���Nr��5*�]ù{A(N6��ZX�͎����^���C�?o�U:��U!���ǵ4��E
@-�����z-�y��}���ĳu��N��S��Ƥھ�9���5�T��o�0ܭ�w�oqm�
�lM;�cqK��i��AHa-AQn��&�S;��H?��i��dK,�&R,M�� *d���x�y�5{�O�>�K�p��c�}:�,!��' �wY�%?��7[d�ÂY��բ��G�����Y��o[��DC��$T�f)̡��a�	E|����b񼈘?�G`:'6�Q���a1i�d�E��8*@�`_{�,�!KjH~�L������;m���<7��	�0�3�o4Ч,��u��s{����Ƙ5�¢���M�}Q�*4D�-'�4w]��)�ED������+��r�D�!��${�klT�u���q;�o��ˆ6���%���G���*u�9=>��a����@�"�8����a=g �l��~R+�ּ���nU!�'��v�6-�EA�����oIX���n����}� QXM�َs��od�h��=���?�o�J�����i=�6�kӒz�#:����GI�W^�so)�����Z|Nir�pj8V�fam_5	<�y�n��qY�6�VѼ�ԠN�xo�Q\:9}��^�%�����+ڍP�o�����40a�5�}��7)���?���7��������]gmD��-�v�N�)9^�/��hfdCӖ)���r�+�Ԥwۢ�[p�؀��;,��Zہ�6q #5��ğ�4o�K� k!��$�6���V�K������6e^�7��"�����%+k�VN!-�*S��� �� �Sr|�MXGT��w�4�����O̲·�<6!u&S�k����x�~��]���'R����>��Tه�8WLa��O�*�,!�o����㰫K�e*�(����/8=.^�!��f�"��$ޒ�c��ڧ�Aa w�.̞D �1�A��u���`ԇ����������9p� P'��w���f�LQ���&��i.���;������-Q��

��"���������+�^&��!�*֏��.n�# ��=(�ZΧ��(ا��q
����X�{}�W�A�Evr��٩p�'��g鮹�|�Z^.��P�����9dgd��))Z��/v����0�� ��i��@aR����$�Ƕ+���*��^L}�f	쵴F����T1� S�k�x�J}�i�zB(?�����A*�1I���4��Lw�Hn�R�5��gͼ�=�b*Ǽ�+�N\�nj5���b���[��E��R�\H4�V�N%�7r��3|�B�hB\��M[m!��- ��P4B���P�����~mTܡc�Yz1F��{��MJ��8�*(�ʃ�����_�����(��l�Ejq��E@�?��\��^3[���-j7x��1��F��/ ;��-─olJ�-il�|~����#�����e5��,�9"�C�h�+U���y_�����7���j#��{��j�4�'IZ��1���&T꼐��R�P��QU�a�a�si��Ԋ[��̎,�Ԅ/G
�I~�������1���dX����$���}r�4�r���L�c-��nV�{1�+iQ�Tl�*�ƦU���U�����\�,LY���7]�,�~�c0>������N������7�#�Q��/�ˌO}�r��t�ر��������*��XW'�E��u�,D���Q:�ih�՘��p2狛m��N�2��AaU�ikk��1W��=VZo��i�{�.�e?ӹ�*�aO+�����Pb�i�׆�fr�x�n#��Ӑ�]Ʃ0	і1I�V�R5��nh��il��>���¼=^� .-y��Ȗ�7I���1Hmj\�Gn�b~ ߏ����#p��� '�>�=�J/ה9�-egh�:7����ɍ7��?=��G����X�,�2�!t'��NBB#ƙ}OX����-,���^P@�9]�hN��2I^̥Fmx~��9ݭ�<�8�;^_d1�4m4!�r�/<��ҏ��� �M@��Ҥg� �)�D[��	y����#��z���G���lPH������8f�r��v�sO44��f��S��0��f�L�%��e����m���"�L����򜈪eP�k�6�껜,����+�6�a���q�2;�ʡ��w��V(҂R�	�w��P=��\K�s��yy��^!�KK��g֮���ΪР���E�(Y���9Ou{t�8&a%i��b(�� �<�ބ�m~F���ia_qN9�\}�IC,0j���.C�Jǌ_V�@�oYo��.3�!�r�/[�c�q������F�`�������Q�BNH#�c�,p�0;t�>�=
S,�]��[#HoS>����҃t�����X ?��l��2&��x�\�S�Y��u "$>�/eÞol��UFwh��.���Tj�Ş�*uVZ�k�pv'���s�T�ϥ`�������8��K2OG_FW
�W�O�;����Ń��۳3�4�h|V��)"Ⱦ�iv�8�@{vz�gf��������[$X��\��&���д^OX�Wb�f�-{�v�S�o�G{2`�b)��(+��	ЛE��}��p�WG"�������M���Ia�n�����K��oA�F�a�oo���
E�n��2Z̊���
<���@���J��L�������y�aV���IR��F�����lױZ?g�����MM�U�}���
7z݃G�D��(�iֲ���-�,l�8���kQ��\��E�V�ŜI��@E�װ��C���0f�2�[�0f~���sϹ�&Y����R�T�-�y��S���G��_IX���h�F�l�8���P�F�B��6�".I������=��R��H�!_�F�`I�D�Ԭ*~8�\�mZ���ߑz�=�k���+ ��Xp�T6�З%5���<�ʠl���S���3��v�΢G^����n�	������ a�g?�w�����W�Q�M���y�����V��*��W���S�`�c��N�VY,�\�4��3�N��m�p.�R"�Bb�i�s��-�1�Lw5oI�|۳��Y�2��=̛b;��}�`��C��yŊ	8%�H���-�B7m�!�#�v�!P��{�p�P����S*�N��!Y��9��k�~P3;���y�hM�ɏ���]*�����`ۼ���@Zy9Ǫ�� f��T�U����|�N~�'�x+�~�G���D�&i��Æ�cUv�!K���3;ڿ�Xs/��Y�i��w�<����&��P�@o:k8as��V>&�J�yn�����������t�	�`{K�Y����s	�����b�>���F/d#pJc@�1�#����.¯ǰJD�	���;ut?e�};|��	�S�+g.��M8sYɺ����Ⲷ�T������Dӓ5a�_�024Ǖ��>�q�@���*6��p�g�@�y̗�8~;����f��
O���ѣ��ǡD`O|/>?�O
���z�F��ۨ �'"�<�k�O�i*��r�O2�wP� ����3lq����u�'f��z�Rg�eI(5`dٙ�If�I�2E-
�Fą�ǁ��b��s�K���?t���z������������A�d�ҭn�
Ix��u�#���$3�[
 �m*ձ�aƊ�R��JLǸ2�2�����ӫl�;��G�� $U�V�1��K���c9�A�sEr��T	�$�t������X�U����6?�}���o�����᫕ΔA�e��1�ZIn,G��}/s`�ܗ�"ș���t(��_��A��zE(���Z$�B":�`�����ݬ#��vY�04�6~c���;Y_�ҕ������/J��j������U�>`��ͣq~�[
�4f9�w�y�� ��M���;M5߱�!�#����b�B2���������{<�p��C�}��[����&Lo�Y���f�)��QN2�_�Wi��5�#���&_� \7Z���wj��}&�
��U�4�IPN�*�_�*3�w��n{p����G��@̯������4ڴ���҈ %X���?@+r��'4�(#���������|���v�pg]��O9��6����};ʳ������uף
p:�	�N���4�Y� ��k_l�?���Yu�Q{�M������\�l���k�1�� ����$����԰ɇ�h��@P�9��|�������� ,ŀ��f"���N�'��	�'?�Q7��"�B0������!�ݐ҅g��Ky������
([դi͂�uv�w`�
S_���.0iⳄ?��r0�CƤ4C����֝+��(�P���(t��Fs�S��<�w���҆�1o����\��1�2Qt��G��H�b9~4uCkWR&�� :m��AWX�s�ۯ`T�p�q�@�f�w�uXܶ)/:�F#~�스��U�e�\��>&l>V����+�&}��@�ʺ���pz����D�&�ۭ��.��͠��)�,�	�'�+��� �V��V �w	���BN��s�������jFQ'�Ë�l�o���,�g���>��V�2���<���5d������P�:�D)�I�l����:���-}`פ�Ȉ獴;Kzب�茶sr����6Pϭ_�dSCy��B� ��W�ܷ�R�l�����H����'�|@�@�i���2�s6b��W���G�i�`
�d:|�.n�u���71�L���=���4�N�l\@��&),�~��x�閖G��S�W�6�=��2N��EW�jv��!=�@Р�r�Ē&n����y���ּ/Μ�v)�DM�7�WP�9��8ؔ��jN)�1$���D��ڤ����<?����%�l	F!�Y�'c���DY(�楟7 �'�X4�	p,����<���E���}U��Ϛ���g��e>�p��5ԯ�dTYw�����U}��`RAU^}Og^Pr�˴W���
�d��D�*Xu��e�>}��2��j�.*_��Z+���|O=� CB[%�{��������B ϼ��<�p%�+5�<$�-Q�V���t�ҧ�y��G��K�����ɭ��4U��Nى����<a���������ê�liX~ 'u��`snf�̈������^��L���8�bxنE���(����� �d��|����n�;e��<�Z��̷��z�#O�ӵ���{��]w���2�D!l�b� ���T��+��؅70t;O���x}�K2�&�8� ���M@xh�y�wO�U�C��Ymn�K�|\�è���Zw��r�PK�8v}.=��6��yY@"������oh��*�(/����@c#h��-�bt5'�u�7�^�f��su�)E&�+�(,-�6�i��ݡ=�ٺ��g����rT��k��iu��D9*�<�@*)8��	�J '�Dx��u������x�]S��J
`�-�İhS$��o@(U��NxmE,��&�OUR���(�&���aږT�K�L{��}ɵ=,==]��4��n�3<��lu˻��/ɹ�����'T��I�	i�,���"�%K<L�?�8%+m�画���p*|5���q6��/�I ?{u��U߲6�� ��d9 �H�=ͮ�_-6_D%�җ��(��7<'�*ܽ����e��&�È{{��fX��X����28��@Ё��B�,5� `�53~!�M�������G�{�|��8�@��m�a���[i䬬��+r�P0S\�%u��,:�A�q��J�T��Y��Va�<���� E3f����<��� �7�y�|�T?D��l1j��z��;#$����o^�h8��r�������MaF���aB{��!�Tp-ᴗ�h�����ZZɢ�ޜ�.�1{ ��{8���t��#��4�#��٩�;&8R�?}�[�:ȡ_l������s�6�l@�f�3(��oo�^*��d�|:��Y���*Z@��'��2j7�HK����O��n�`l��K�[�c%�"Ώ��A������_�p�.�&�m��O���i��ο<*�+�n<5E9���xShO�B�s�S�.���Ի.me��^�P���dN�'�&W��<��{�݌���]��$�&_�݅�_���z�!���P4QBĄ5߇Z"mH^�҃D�Hz���6��k���������rD�|��G���C��;�_��]Y�˿������z�<�
/k�JڼHY����@�/�!��� v��b�W`st����f^0�����~�����|�P���+�D��|��Y���8#���xj�`�5���(F�W�1Ӽ'�Av�l���TO�贇ϟө ��v�,tM2۴�{Rq������m(��k�E��;!f���CÞ�U �/kD����aW�����Y�Ⱥ��^�v��>�W<�gG���7��0e��$��#Fɘ�O��.���ɟ�+�W�Ϫ�;(��t\�<����T��ᄻ��Z���]^pʗ���a���(��Z\>0I��Aj�jQ�G�p���O�";��0��h"3�x'���~0tb�/H�ڬ��A��Ɗ�͇Q�����+V�\f��[����2�o��`�SU�����*���#1�60v��d!pGvWr��O��#����/d����ą��+�6_�&�f���Ի�X@�ox(y��w>}3��㠲�eb�8�M4J��(���n"D�1{êA'u�:����V�#��5�q^���>9C��7uu����j���0�̽<�c]Y}�vG��%}�'s?�[Oy�0�'��r���Uztx�b�^���)��){����5/q�4�2Iռ�����N�M�uo��������R|O`XW�g�xD����i���T�E+�U��`��h�����B��XB�LEl\��$�yJ.q�F�"��F������$�d���+,�KM��'�\�d(�_�j	�K��Y䙔�r:����e�+c�� $��C��
�!,n��N?���ߠ�ٙ���ݤ�}=9ےX{"fQ+�%��I̮���Q�7�inx~ ��jҙ]C	xk-uk�!~�%$�G/,Dy����#Y�'咎
�S`u� �a�E��C�ew�>c�t�]68�32M�_S�;5��=��x����9j��T���#���^^�]j��KY�Jst�@�����jg���	d}�»���m!53�#rwT�Q+N����C�� ���O>
U!�ԅ����Qw^�m_n�l���Ӡӷ�#
b��ϲ�F��z]���k�l��Ik`o�s�:�=�s�ԣ��G7�^��8�6�Llĉ��6껬[���BI������Lm��z�\���3�d�]�h*H ��k�����U�w���c�1��_=�.@.�������t�(���ú����˒���SȽ)���҇;X�֓��K�0��1� y�vNn:��-��&���M� ���jǙs�w����0�G�X�l��HW.~�~�g�Z��S��q��������k�B�H�?�z��ݯ��!N���T(5*�8c��^9p��	��%Ԫ�
��S���^���8�#:҃6���wK�.5f�V�:5��)��lY!�q�s�� �|�\�p6@�]�5sI݊T;#���Њ��C�����ԍ��X�8�z"IT�<�v9��Q����I9Z�LT��d�v�^;t����[��0M�{C�ML?��G4���]!j�QZ#��u4��6| L��_�ggi?�3��=��9�n��'�	�٥�H�_��Nը�K���S
�P2�i��H�v!�ł��Rc�����߆�Y�6���O�T~dYbv�}�Z}BWY�k���F�qf�������d}w�X�>T���P�_K�������E�LO������%����>Fd��oj*��$��(�VT;���v=�K�#S4]K$	H��E3�h�,����t2��)���=ElhuY��a���Y�Ґh�x�kH�x��ަ0�����zM�H��)�ڋ�@����9�7���[��D�PJ��|��늭5l<�llҐi b0N�d��7ր��c��Z�iܳ��TF��}�<*p��dr����
lh\W�%>)4� �k��+��b���Ke� a��cm�[,Ep�&qї��؅w�=4a�)�#i������כ���M�/�y3�,2|�����qR�c�/ޗ�F��YSF�BÇ�}����t��6�h���+�}P�s�ǀ4Lky�v��ߌ�m.]~F|�׊��$E��3%���;1
j@g����f�V28�v��J�ۤν0gQ��	��9�aqڻ*��a?$ �`����E�cf�g�[�ۖ�Ç*&��^q�:�@�Ju)�4wx���H���Sw�<]��%����-[a�O~p��d,w�2�����=�Z��` =�{�dړr�	��,	q�*)U���/#�� ��8};�F3���E����T���4�'D�2���3��eM ���PnL�8�x��)�\���>�yX*ͯ�/��<�4�P ������p1[|�+9i��!�z*�!��}}��ED�5BB=�!��S+Ff���>��bR�w��x(ے/s1�j�uo~��W����LZ��y�s�.�*���嚓&]�e��\G�A��u�`��dKEm��h�j��j����ҤG�_c��op���E����V�xW��ILMy9xT	`@ݽ�jJ����x�Z�
���8��FW�T�4W�	[���t�΋��ޔ��vbr2�C��CnI�j&=߁��������|z�N{6�;���$�)���J+�\\�!��*���4O&Nj~��%�sX_N?�VV��}uaB�s��04���˼��RX�!��%�Yw"�f�4Ew�n���3 F����g���!��Mr����iR]����ocg1��D�����Q�ȥŃ��*�?�HwM�*��:�V�H�r��3��)�Hl�}:�(�.�-'�D�Q�݁Z�Z�Uf��mͰ�%�8�_O���Uf�M��zQP�3ž�I��Z�
���� Z���3�[����+���-�З�t��������w���a��O�W��?�E�]��a�܀m�$ߙ�q�B$���aq����o?Ε:�2ȕy�y�e�l��-��y�H����F���:�<\�S�u�8�M.�|E�z�I�7Mv�xe�jz`�S��;����YQ��x��8 g�Y��.��� Ǖ�����<����qh��dw.�L�����㿑����S��dݡ6�(�)�dL?5�5^p>�u%�P �T&S��@�΍�cp����P�sN�}أG�	Y�!��@ʒةH-3k.�զ�6q�%�M�����D8E�]���,��R��-�F&OPZ_���U�U�����oT��3S!�?�{�ߚp!,fih���q�A�l��ZKQ#?�_U�W��Ԥ+q���$��Kz��D�)���������o�F-�Iv�`B��ӌ.�b6�P>k�_-l��"'(hU�bzvb�1b�#Ҡ�Q�l�l�/ߡ�P��g��"��$G�v��\*.@m���OV]z�#�ɤ�3w���^��H���l��<�y"<�~az�Q�t���`b���ğ6V,�����V����u�8!��7<�lr�0���<+;q7�/�D����XP�`ao��$t9���.��ޤ�u�����Q|!�h��>����E�S]֨��t���Ek裄�OW��.<��wXD���u��@��*� R�l�#���PTb>�"��� ��6�P�X�'A���(a��]$�V��{AV=OY��6�".iK��!����[����PP����N�0����n:�^�j�F7��ޤ���}���r�mƑ|[NW�V�b�ɠ������K�d����?�}���3�֝qM�Q��,Z���Xy!v��*m{�R��u&��?E#�9j:뛹u�l�O���2�4���1k�����#�D��im��廨R5�S�Ttp5edRx���zLq���u�@�0����]ᭇ,V6YeZ�U=Do��Y�y�C�z�4�#E`b~�Z!b$\/ۑh�}��>6�4q��W�-P��e'�� Ӧ�BAdY�:���GsK��V�F�jx*����𒕡�JhV�)S��h����2|_|�۞^���a�=tx�~m�t}9u�犔����V0Ü�C.�$*� ���Bu	����V̺2A�K3Q�zF"6V���{��^m3��E,�d{���3]i�|wlQ�oL��wO�n�����Sԋ�D���o�?	�Xr�\�3�,�B��;ߕ��"��u��k�q��v���5CW
�)�C��xb�t,}�\�����eGؕ�T��0�	�Vf��	;������rC[gZNL�W�PYGJ|�A��n:5�K�����x��&<Q�6�����T�͊�8�\�Bo��Ð��)20P�f��e�J}d��7N�9+�<G�]�~����+u��A���W71K�S#�"��>�P'̜��3��g����F�M8�a�Z���T�(Z�����Z����I4-��>�Km� e�lt����ީ�Ħ�<]c��������+qw��B�I�i�F��V�1������ޣ�4�89Ub���hcc��E��V��&ehz+�Gt�D1gO���s��h/C���l���~xn��%�h�-)�;߬�9%ˣ�"+c��<<���b).�N�����Y����Q���n�c6d~Tb-�����,�핫�\0�a��ԯ�ݣ�ӷd\�Ҕc¥w^���LXB�f��É;Od�'�v#⟖�6`�ha�{6�h��uOs�r��D���ȒFW����V���"4��<^�;kC����N3�r �JlB�R�V7���A�}��vG�h�b:So�;�f������-���05������� "���w�����D�r��m�H�����dv�bs��?g��+�?�e ��S��'=xҹO�_�_(V̴W��H��XIFU�k���0�wG6Ǩ���۟���xC0���dcj�8���]�`4%�����WH7lTe��� �j��5U$�9���w��q6�;;$����˫��x�P�w��Y��C[&��Rl�V`=�d�~+���>c��C���e�@@�g��A!�^j�'C^�
r��6��H�ʿ�\�	���o�0���������{���rw���u�-B�X��W���?���k��ŖS����5YwY����J�MK���.m\xy�གྷ���e>%:��ᝮ+��J�3{j�q�ԳVB?JI����w3��g|��ݠ���I)^��R6�2&B�t]�w^,���O��M�l��%ߥԶe�`�5�DsX�žc1�S���
8�&�Kn<*l�+P�P\��iqwWp�����݌#'%���m��9��ǌȈ���|��Y��5�������mLo��C��dE�IU9��������li�ϓE�������-�]���4�O���3�����2ꫥ��L:�?���5@1O[�� W����Y�D�I����#��[���rݟC���}��TMd�i8S#�o`��$#�J���a�/���6�0f��~��)���~�㵙.mT����7ܠ�gA��Y9��y�e�Emv�<�7�$ �+|7���4SV����2�ww�;(�1X�{�er+�M���r�xi��T�����#d�X`x�.�����ƥy���j�0j���{ �J��s%���}��d_����L`W=&��B�֢��8h@��ף윣������]�zI7q����a����㰺Kʱ�=a!^���\	�����n_�7'��9�.��eW�A���u���>���P=xU0���'p�cs�@����nCr�iS��Yف���E�X��`P���8۔�pf�b����΁���k�������0cm�`���V��)��E�P�p�#a��Ǟ�����_3�f�������}CQ3�Y  �`WL7���q6����9��2��V��u���#��ڠ��B�<dt��x��U�t���7
��||��6��*G?�!��!v�j��Q��i�')���"S��B:�lۧ8�N�Q0��@gM2�=e�>�g��.������>�V�9����b=�e�����{����,"��$*��]�	���6��~����r�2fJ@���#Ι�P��*I(�Y\��{sV�=�/�����.�dZER�׏�χ���y6��j�[R�!��x��m���F+{��c�ȋ�a�t���>��v����]�H-FU�	z�@ֽדu��x/��M�Ԭ��ly$���xk���}�F�o�S�m��rx�W�`\n;/t�]��[��i���/�~�gie�?�eo�J��͉��0P\\�(a���V�z 1<�5^_��})�:[�v�,��:�Vs�'7���~���z��$6�t:�M��c�����fc�@�g���~��V�P�s=�-�v�M�����t"8��D;�D0�7�%��7z��������B{Y�.whkW�t5i�=]F�8�wۏ���k'����YJ�H!�z�,l!�7���D�����h�˳z��	C��[Q���U�RM�C=�hq౴��7�����%�ɾK06<�]�[�(<r�w�_�^�qћ;�&�S8�ID��w9
��$�)�Gȸ:{%5��	R=���TdN����SI�Cd�;#�J�'=��\��K���>�cJh<Opwbom����t�{�\;0VRtF��)x�hr���BI`^y��B�r�9�~^�m�n+�m�ȑs2�u���A����'���'�7Sfͱ���8�ې��ch0��|W�5�7�����c0�e3�.w�x��0.�����A���xQtT�V����8l��l1y�r�;��K�.�Į}���'a�9��ސ�w�"����֧R8�iG��CZz�[и��Y����S Y�{J��v��j���\���RE~+�'�ZȰ�1uj�l1����:��ȑ%�GT�uJb%|t�(!��i�Y�v���Np�������E?
�p�a3X�����B[�K��:+~p�����0�
s�"�0�$�I��R�姼���#N�e�sv��Y�,aY&��l��i��`!�5�A�jH �(�>5v��:���0�}���܉��4fQ�-D5y*�,�m\���[l�����@,������=��~�K7ߘ-�Z�E� Ϯ�)�ۡxs�4�Ns B�NBdqC���ABUg��_ p�M�3bKՃ���͂_���2��� OAM^��<ȵS�B��.U������J#F���Ll�:XZ{��h�T����]f�+�2#r�J8z��lVig<��@�b���ȓ���u�P8�.�����[���4~������9�B��a�^�|^�K�^���Law ��[���:�KKKD�Es���at�*�b�%��$�l��wzi5�Ǫ(�%a5�/'+B��;�#�J������o�՟��Y�'0G��L�%!I�C�����
��:��o������|ٞ	�k_Ͼ[�zP`(J�bm�����.�rƷյ�w���6������m`�i��ưZ�>��P��lc��'��;�P<j�5e���*˶	�������H+��w�⦏�w�9.0��ε������ZŰ89�d����B�@c�퀴 kK��'����K�L��pH��{��O��` ��ȋ��~<�����������!��LSg�~����L��&��ءL�B�Jz��F�:�����e�y�C}�&����@���hqD$a�;lJ(}��.`E�>`<�8��'��7��N|�[��.�ͼ�"	3�9c�G�3>����lf��N-X�\�/Ң%[�K�R�����t�Tj��&Qe���������f'_��IFm��4�LK9���� �y��η᠟G��wJ'v�wZ0�g��k{">�nh�S��|�G��˜+|�������Z� �I`@;�$$�WJ�M2G��o�H��>Ĭ��44Sf߸A�
*��OZA޽n_KG����Q�Tk����%�	1���͓G����DDkU��R1L0D��Hh�FD�F����[�ؤ��C�f�	
B��0�"G����d'3����=�xͬ�y�"�=k��a�IrP�C^��V*�zxZ�����`��b��dH-ѶB�IO���s��w�5&��m�{�� ��[�5�;>�י�e(Q+YN���ZtG���*?#4��5�LxAQtf��������3{%t
>ץ|TLA�Q�� ���s=7\��=�V��S�Wk?��h�")L�"��S�"??���
5���{�f>�=�X�g�?ʚU�Q�Vir����� Ci ?Z����rlK ^����*%  1L��X��̢�8¶���/b�x#��
!��t�_�]�l��YI�n��B�P�^��;��P�}}�'��;N*!��}��u���,4�K$��G���L�t�#o�]'�C�Z�ӈ�����.�����@N�`�+�O�>xU���{�AN�Q��D���jQ@=�U��&e�
�>�[~K(��>O�D�K����	���t&���J�6`ɶ����?Js4(m��4���U�nY��0C�4{[�Z-MA��eup�2}161\릔��L<}L�����i��Ѫ^{߲d{����V��$X4
�e1��0f�}�͇�v��,��ZV�I��[/�ԭY�Y��"c*�5[iM��m�|�r���?�Q��m���Rq�[�X=�\Q[�K��$��=��^b�𭄚 ��1�����B�Sd���>C��NX&_e�����/t��y�f@b���s�#n/���J\��.�XG�Ŧ��%TC�D?���m���s�$������4Vi#P
�L��rs1z�H����^吿���\;T!a�\r�"�Yz����Oj�Л3+��� P�z[��\�L�O�hh��BFtXZH-:�M�~���%�<�Vܽ���|Ws�lb��:@���,�Uc���E��	�Z]I_GY�]���N~q{ ����ߚP��x�fHY�_<H���tYb�귄2$̀3J�������S����;�o�}J�r�\��k���� �A��nW.L-3ԍZM�q��\۲�sd�~�P��f�[�&�S�K���˸��R8Z��Ӥ=ݵlV����׌ޘ�8��8vw�ŞdZCEe4�4���y�S�����-i�/��se�d�Mu�(+��Ƭ�a�V�j&�v
�E���[�0֜�-����6�\o�f������h:v������N�����������N�W�\];�1�T}�3
�MX��^��e���y��� _0���g�ۮ*���������mP�C�a>�a������r`z[�TC܋���&�'��c�CC�����ƀ��I^�٢y��x�Up�&�{
_jk%$竐>B&�!Y,5ݨ�J�v���!Ih��
~
>@^|&�岑���*.�G�P�-�׸�� �<������GԒ0��j
k�-!rs�<���NW��I��֋��΂�4f��pB�@P.mfO�ɐ�J�m���Y���	�F�n�gPD� �O��pbŜ�!���+V��3H�����Su��q�G�]]nQhk6��2FX�c^<���F�8�1�]8&	�ߢ�!��[jb�E@�k-���}n�����x�N#��x%�c�V�޺Q��K�b���{4j�g'[��t$+`#�3����V6ھ�);�YN�z�/�a�5Ücdo�=;R����K������h
/���-�j�^���>j@ٮ#J��t�XC��qi��vB���i���N���i���xd�
3γ��,���)��\YG�>Y%j�F��jp$�����.b �}��³�U7�1��-ע���eE����$M��}x�#��drdPF����z��mDO�WeE$�R�
q�wo�NQ=��1�o�
?R=�2ո�;=�`9���`����?P���l�~R�p�۲�2�qE��4�?O��4~���C�y�2>�A��v�����9$ʰ'����������M}.�in�7!��0yVLȤ-�*�M��(�IG�xg�2H7�̏ܬn��籢��}�ֶW�^����t!uo`/~u���g�z0}�8�@r��]�ߐ`�l��x={��Ddu�=۟snƢ5J &���}Ө��,�R�װw�.C�u�_���lǫUg+$��2@/��A뺴�s�D~����gk/�wp���;Zǉ�h�{��r�c��&/ؙ�=j��{��^����aD)�w�m�a��������X\���Ak��!v�N;��A6���T{�q��R��S7��*�)Uk8t�hg�|��Ǒs3H��K�qO�ps�P��i�c�U{�����͗�r���(�eO_(��!S���/�i�J	�1��-�sMX������w� ䷛���Q�x)8�L\��V��rw�V�˼�: IfΠ
//=	���
[@/pb02��~C߉7�IM�J�rt�Ώ����Z��9Y� �sN��3o������lχ63����@CO^ti�j����#�����ml�@8_wӼ��š����T�n�[#�[Rw�z��Gn�Vgb���Ӷo�[D�J-H�`�C�%7�Q�vE�W��0h�BQٟҀ�Fľ���Gb�J�I�I:�<^t� �x5�}��V]�J���I8���8�1$5Z��w�C��F�͑^HSR_p���V6�P���jÀ������M��*�vp��)��'Д~�2Z
�������T,A���&�6 ���$��^X�K�[ǟaDD(��/*;_��>�(��wj�|�ze7khx�#Z�VԂ�
V/���5���(�j$��4r��e��X�����,=�l�h�Z'����*:0j���f+?E5�F��!S��;}�rd��&��{��M�-���u�贐ݸ���5&s�ƍ�0��و�6�T 
�O������D�OHԔ^b�d#�N��j��C"�ehFm#>�P�٢+��1��T��ޮ����8d �m�i��:5��+���qs����/�9���b8�D V���$\�C�#,1	ז�������f^��Q�!�̣׾s�z�&���sA�~p��F۩�ڡ)�$�������l3��g�$�0�8B5y�b���~+�o��ų��0��vN�.6�Xк-�+8��_�-���Z&���u�Q���ϑ�HvІ�q��6�-������p�j��;���+��.ܞn�6��.@�ѽa{�#F3ځ�#R�u����9k�?L/���{%j��v����P�F,>��A[�N�u�y>h�C�G��*����f�����߸�����o��I�+����c2D�^[<�~'��1$AZ�w��ρ�7�������/W�z���N*k�灾G���F�uNL�rB�T�]�?/\�,d�9����2�X P���_C;��ˏ�����Q4䛷�~����aN���z�^�R�,�ǚ��4U�@{��&��˶j��tZ�=�jmH�vp�|���>e��[�H~��K^�0 "��;7�G��C}����*އz�����K[��'5���p��z�������햍�g1�@��׏r��s���X[;�2�R�(���(��U�U�Ð���ɱo��[{�W����t�����oq�����ޗ���K�p���������
���j"��7��s�V�c�I�Ea�.��ӥ��i�(�j�c��ik�~�ߜ�xS*�-d+�֞���-�-8tT)��i�d.�c<V�OL_�Jfd���5��'��\Cpd3�N8���ь�s��8]�֏����cl���A��|C�����C��|T�X�=�}�.�/��/�۫����Q�"Q���ru�3�#����V� ��]W�
��&�H�����	���)��/YʠPY����[��Cj��K<0���f>����ѷ)��bc���A�U��lj�0�D�~dl��[y�B��IZ8�JR	n���[*Ȕޫ�)?�)�C�j*�ecX*��HߙR��|�=̵���K�8"9|IeX���MFGu��VR�ޣ���pC{`��Ƨ}�ٍ.�|�6�P"[1'j�G��������2�-��X��"�O���@�<�9]\G�9o^ˉ���W��B�0�\�)���@oDo�8.w��8��w'A�EAvwaE�����P�Po�A�&-�o�<H�#�]�ɗEl��p�e�<%�{�Vl�R䰻E7�Hd�M�f_�@�}Y�9I0Y�
'_i_�@K�_� ���M�![3�"Hek\��/sN���7zb�i�g��wl= �K�������8�
�K)ql�'q��&E�z�Ga��R~u�oEL*u�snf�]zB)/0�r�� fM���bF%��ͻH��ɩ�V7�/��[L[8gPD:o['KdVj�h�`�ԕ��ȵY�a�
M)�^�#3L�tN�H`y����A��a��|�_�l�G��MifqjX,D?���/`���A���C΀{5R��p�"�"�B�������̈́���Op�6�F$����x���uɼI>�6�ܧ�����9�KFYM�j�$�1��\[YtS��J�e�������Ou��q袨F��pw��������.�ٌIg������w��f�2��Wq
?e : ��xI��|�!pE3^�q�}�AA�v�4�z�d�����Ay��AZDZ'�65��[��[^9��6	f��U�w~��W�.C�͹��k*��.�]�Z�$
�$[ �Y�����7�M�_���t���@1�����ѕ��y(��8�y|�M���F��?o"������sE�e��9�`=��zlQ�h4�`g���4A��v�n��i
��2�x�I5�����\�`��+ג��?<I%�Q�~P7Y�]Qf:si�O�Yr�N�y�.P����`k�����G�R����)Is=�7�ҙC�Xu �������w���e�%��#9KUp��C�$$�x��w)���7��<F}@����u]Q�뱤�,[�@��N�O�@����˯Ѥ�A.�F=5�#�y{E�V쫜�*����̉�L6�D7�n�^������Vj}�oZ�I��0�n]T�o����!$�2�zi���FDt��??�N�*�_�W�a
�O�N�<�u�|8;���/s,5qI���
P��{�6t��x�@�����Z�ce�������C�s�Ƙ�o�U�,�h85�W�m���,��ac#��V�i���p�%5�/� �a�oݍ�RQK�=��%͛���Ѻ����Q�d�zG�+�9��q`B��q�u�y,U��xA_,Hkp�oLɧ=�m)���6��Њ��N���Q�s����|��X�|+.�X��ׇ���N����.6'�za�2nR��SC��b���>A'c4��j6:���β}���M�1�y�E0�j�9�_�6�{_5���8�w�ȝ���$��������ȿH��9l�e�O�2�鬄��﫛&�L�N&�J� �W1U��he��F+�u�Z���M�AVן��Vӆ+����Q�W=4���)]��w4E�W��d�C�t L�!{�Ffz���W)`?�胁�ν��;2/�d'�� x/3s�	�@����y�������o����1�v�	�Rf�yEl{������W�Ǒht8� bݿ����!�6.i݂;��Vm{H(�}���s󩧨�h�y���\W�pT�e�S�x���(դ��H'�1�ԙbPQ#�MÎ����0���.�UbIW��+�[f��ձ a5gR���4^`��%��<Y�T�Ӕ��oj�]��h�ZR�á��[��K�xI��*b��4�)��z��|Ѻ�ww�wt��*!-��aA ��S>4��w5K�0~�B��6�g���4K�s��4�Ew�+@N���l�o9U���v�qd��:l��Ag�Б�� �쐳���IH|>�^�X�I�N����Ix�7���v�7
��ǲ��Wn?TQg�����y@�K�G�װ�|o�y.=l
�4����,z��*M1��~�#ęI6>���"�J>V�ʕ}��N�6�T�������,3a�G�?�j�z���b��s�h;��=��%����ӠMI�c�:��;SV��Cbh3r���/
��ST�?��G%�7)�a�1"wA�Ӷ�^b���u�dK��:�25�¯axs�͸��יمԥ��R�&vA����Q`��7W����7-�o�M�w�̀�����? `9g��{�>0K��6�W��]��X�U�a�>�vn��A \��Tى�:za��V4����w)Lt:8/�z.���X�V��[Ȑ�3P�VZ�h+M�ٟ�b���l�\�D�]�	��՞�ㆻ���fx��fA<�p�*��.˖bݶ}>���#%�g�r�QƏR{����w�a�z��32�w�0w ��	n���oe>�IzmH�F�hi�V��"'/�E�yC���P%�D����b�͙a��*GK���6)aX���c�[���	٬�j���\��3Nx��&o�Y�3���FN�n��� Mh3��&��΁5ɂ����-E'�A^�w,k*��X��4�!�<X�F�c0h��-L���fj]�e`�D���}�˂�p�%n�3`�&ۉX��"p�?.{�����}�#�pӠ��?cM[����p Z<�(�!Y#�8.��_ Gq`�y�SQM����<��O=�e�xv��q# {��R��"���DV��򺌴���|[���	2��ȪÉ��kOJȮ0��J�[	�ج?M�#�@t蒦?����h�wՠ���A	z5�A�[6��
f�
~3Uv��o5�ĩ�'2�x\R�`�[�VT�y�� �d+.6�������z�F@�0�cW�k
��oyeT�xc��q�l�[��~�x�Y���x�b��۫���cV4��gO������%O���`��e ��>�J�[����M%�"�|�%��q�_ü�o�X�c>�V����JY�]#b�S��\AZ�.�a�4��3��:=E���t��Qॲ�!�-��g��'�z@)=��A��H��A���������n��V<��M+�qӺ���_v������79��^�����q��t랫)<ԡZp��i:�A�h��3����K���=��J���4�`�~��7Sҏ_����u�*+���d@oݷV/r=G�����4P��Ff�J$��Qa��/r����d��[#+���5��v�K�-��Ki��6���h���.ծ�!���hI����������C�(#�=��M�B�=W �0C��ONC����Dr#��Ts����w�<d�&Ţ?K��x�g�3�Իn���R�i�t�ۘ���:#�;2C�k�f����/ᛐ�qH'���9li��Du¸�A�Nڞ|�p4�}�������d�5WQ���	���m֩n[��"���Xڰ�~�s�l�c���a��a7���R+U%_�|Q15�L�S+cQ��l�+�"�KwLE,�xYo.&�QGW> +b\��z��e S��K�կ�Fl�u�#��n�7W�dQs��@�B/�k+f���%&I ���t��ti��X⯙��6�<`�?�����tp��Z���$�7:�_�$nf]풹%YKٰF+�o����  ��܄�f��wp�+3�7)~�f���� <����F�����Z_�_#nޤ�Ä�>k�������s�j��.��Kf}�~�����#A,���J�§RD���M�r���t�7S&���~D[��o�|_R������%=�\��J��mD7��H=5tQ�qMǔ��&I���f��?l=ąXU��\f{}�y�rвsGW�8�s��8�5(�*n���Ȉg����Oǧ[�h��+BՕx�ƨ�K(#Έo�u=�ҍ	SeB�g,\�� `.��X�4ОS]��g�����z��������	Rƫ��(���3��,��c��P�vi�&e��m���!c�x��������(�]���G�w_\[rŊF	�DU[ ��V��-������RbՔ���K���||�F��=���.���=3�g\���|�Ң���p���X�e�t5����Ȱ�ӆ&d���S˵f�f��lZ�'g�ܧ��)��+�\��޴��nQ��]�N�V�(�b�d���F�n�C�xue�s�y�&������� P����-��oD;�`�(��_��u\�>3���)�@AmH��CJ_�:�h���ҝL�PR>o�����^aN)��	d�w�[�Im���w�_�p=�I��~�[����5��G�d6\/��(��"R�e֢��s�8[�1��8d���>2{'��:]9�v�d~�pp ;�#0B�W}H�1:>^l�7���@_���mq*���ݶ��"��W�B
ߊ��pL�}ti݄�Խ�#���ҟ@v�&ব���6��)!�W��s��������5?q��]�}����{a������I�]��?��ʔ���(/ Ba�(�y`���طr�86�28k�`S�+׮&�� �=�A5�����Z��)�';7�y<>(-����s"Rq�%:�+���u3MΦ�}����p/�!�aX�<.}|�j�ٵz=�5����c�K�"�xz0�#i�3~Ak�AoU<�ӱ�Xm�	>��|�G+��� �o���fۻ9��ǳ�$��IT�53�3-����k$د�#�&%'ű���YQn^�A:�5!!Sv�;5 �-�m�^
E������۳���/"�I
�&�������g����,��d;��͗�y��#�>s�/�#��x���>��>U1I'��e
0>��~�~OF�j��JЗ$�Dr�۶�vN�W!�N���_m��a�C%�-Bx3�!F���%�vrك��Hd�g���nVk��1�~�-�hP��9E����Ѹw�[vREp����H�(esJ˖��9�H�_*	��:mg�t�"��<.+Ty|H�Ǿ��	����*�������ǐ�H=�?7u����U�<� %�|+'w���_zJ>۪�0Β����C��b�s�@O7g��8!�0��2�,�P0��Z2�ȅ�6�k������1�\.�����b��jA�S�6�,f)�O���xs��E�NR�c���]3z�o���@q�B��u+���ju�>����C��Ǘ�Hw9�Ʋ��&-��&�k-����-�ڭ-��z"1�+t 4͆�Bq���?����0*�K���El�~v���hq2��|�����;�nK��{��RJ����WcfؖMYf���x�\�L�O) �X��r�a��z����10�ᆠV�4u�2!P�;�X��3�́wKVy��s��n�����8,�F�+ �b(�oX��Ĥ��󤥰;���ũ����P�a!H���[��P����엿,�l��{��25�)����1ή������q��Lv��-l%��mms*s~mY��X^\P�5(����I�R��W�豝��b���%�����ګĺfQ��
{����מ]i�@!��l�4�DR�O�C4y�'h�,���N�4wF�Eq8R���ϙ�G�&������0�V�|!d�p*K�Dk_�
ߍ�EHt�3JA�r��4Ћ]cط;3���D��/�j�Ub���DV��P� 2k���:u�.���@�b���_�^�9N��.Qk��}8/���Gؘ�X�adJ��R� |̀���~�r�-��|S�I����&<x���b�L����6��j��+��A=���j�6x�.�
;Z8�=v�O/JA�$�rj����.N���M�)nH�ۊ�¸V>&j<��4��b��WE\�y3��� ��2v�e��D�NK�J?�)et�*r��``�� U��s�@)F�lOB�8��/�yƬ/A����ktrN�V~ ���쯷��Y<�F_�^�r
J[�RC�QV�5��al|�u����ڊ�̱��K6Sr�Y4�Xu�vXŌI&2�2�AY-K"���jO��2���:�c'*w����ak��9U&������`��PD����JP3�|��(�(�j�%A�x2��RG\ޭ*�~Y�k(?L�=�7 �܌�vP�Pn��pc�o�������T1�Fp�Ӻ(���N�z�"^�y�>c!ՓNgw�z�\����1��C� �n�v|�"�gˁ��#O\+�DkMj�
����/ �?��Zvo���A��  �u�!)����>Hab�*A� yE]U���^-"vF�1�q�������g��Fd6�$�G��^�'���+14{���&u�q[O�0[DNx$!��r�C�a�*����,�K�ϊ�ݻE�*�1�&��;2�%���-.�F�I��~1�5)]"u��`Ռda�jq,�s'��+��0�aS)�׏E�0:��������3&�	7�ȋx<�?,.�
y�y��1��~0��c�=)Q�N��A��u���]�+��R!�`�6�֨3sK����kH��]V���l�+�ԣ<�W*o��U�0���Ϫ�u�`ٴ�9�%�#���X?AC>�%�o����;���4�{& wW����<�iRLߗ+�'�=F��?�B��$lbe��&���c��sY��w��;�CUҪғB˩	F*��ۻ��V�q{]ڹŦ���Z�<W��9��!����E�@��5��'6)���i������NRył�$�����I��$�^��35=P�e��"���(vB�k�s��l�b~9���\;�1�\��)V��{gjZ(WB��<V�d[ǹ0��,�+iFF����L��>��8iԈ�����vIl��Vrm=�!xXo���/�:wL��ч�hR4��z!3��w�hb�U��b֟h#�e��U�D���cӾJ�zp��	�O�R8ցfǙ�4<�p8va��ub��r(Y^���34
W��a=��<w�ݻ�򚳘��#ߤ6�>㢝s���ԭ����o��"�@�Օz�xv�Ih�J�ū����fK;�rD��=��;��H��/�d��C�9�>ILU^B�;���Y�	�y��?�A�Y���H/S�|���Y�����m2� �u�E����O����v2�G{W2\T9s�l�:�#��Q7
ݭ���A�5_=9���ioQ)D��Hy�?�0<}��L��W(KV�ۓ@��E{�x�L׋���=<��o7���V3鍇i���=q��TC��;|�;�؇�@������ծ4�=���#�p�G�V��؉æ�&i_����%���\Q�5�L�t��^�&\��4ygb�cm>iO��W����9%>�v��C��/���E�X�/�?Όk�7"L�VבL,1�*1�=Iԍ`��5��sL��%�c�4F���ż觋���M�8�6A�.�X
+��p�B</�5�׺��A/�w���Ӕ�ǭ��dD��'�����n�+�:�:�W<,@o)FK7A~��ص�F3o�h�ħO���E��;�]Gz����-{�ێ��o�a�!����߳zr�5��<\��K���DVD�l�m����}�"�Q͗$��[JtD��I'��k�|J�ԩ��.2���3�2$|��,�5qB��߭"�_�m�N��)Wg�?�뇒죥'��~���LL�G�g"�d�?'2�b�H���Rg0̪1uF�&6��9��V�q��h�����/DA����9U@}��$�z�2?EVdՎ<�_���WTC�l�D�����	&�x?����7�:V�~h��а�d9��e��瞖�4�n����r������r���$�J?^�FM縬9]�/Z�_����Ƚ*Y(�h�i���[P�V�&�>#ul_��VӨ�	גJE?���NWX1Q2��|�¸B�b�	��6��TV綊x�7C��-<Ī֓ҥ����'{����|�	 $�=0��&����a��I�ǝ�t��)a� b��l���h�Wl�\�,v�(����$u��W~�� �Oj��0G�88f�@j=��؋���ټ��B-�yc��!�?�k$�lY�<(T���|V%�:Ȱ;Ǿ�
� ��c�Gb������w zw	u�A��D�w���Be@>׷�*ǲ�j
����G/D����}��8�5�:�'�&���+V��1�,L�>|��&�t1'��:�n��986ع�1��0m�L�R����V�*0�h���z���+ui�����#�kI1u9>A-�Ò�ӻ핖^OW+�s�������( ���'�I�ѫ�����0��?�7�{� ~@��8002"����3��{��Z�7��h�N���P(���X\���� ����Y�y�#�%�� W�w��K��8�N��O ���(���/��M1���;J�d@�9@�lWx�`�p\`� {؈���#6�M7rϮ���� ��aS��9]0���P�4���e����#Ve�2�*�N�ԅd_����L[�uh� qL���fh"pr���*N���kg�S ��i�� �3i�_7�I����
�ŜR�a�VωzS��'$X��V6�h%� �(
ə�T�atTYX��i0t��ŕ���|=J$?.��A�O�X�@_&�m�<�q䨴`0�o�.2 KTT*ؘ���PY@�y���5�C��K3�kV�)�c웩N� 3�b������_,��v���9�3O���5 �%���x��l #�Ê����#E^,3��>/�k��Uٵ�ҳ�]�	���r�������v�<��ٲ'�(���5�����L��a�y�� rÐ���˅-<��V�5�j"r{��[�+G����6����k��ųu%�s3�x`�r ��k���Rf�*�FSq��fӕZ��ZS����ޥL�>�?�'%�Nކ��*���B��?��y��h8k����8>�|�{�X�6�'SP;�ӆY�<`�K�>Q���#:Ӡ����zZ�2Pu�B�N��8���Ǽ�AfKEk9��t�J�06lJC�0��<eQa���<_������H�K?�g}�ܘkx�+��=�dVש���6�9!\��Ǵ�7ܾ�'o�A��HL_�e,��2������I�N��w�]�Բ���ǥ �+d�H�!��[B�;����e�DVŠD�'�0�3����N�Va<b��M�'{.ȶ��Q4��m{�HͲ��)U��!�o�~r��8ST�bM�/��-�}U�ju�l���Ї�*����k�>:�kh\����"-�Mر�AxHg
��a"��@7sV��[C��w�Z	@&Qu�����j̐6�t�.�g���6����K�K���X0j/e��(;3C��T�Pu٣Sal}�b��������d��>�.��5
n���%�mq�uTTLi!j)� C��n2���*�����Pl�Y?W�d
Ary���#�a?��(��&h������d�E�����&�������p�XJGA�D������S��.T:����f-����m_3��^oڏ$�������|&�*�7-�������$ɸȢ����ܙ����Qq���/����@`�[m��Xߓא��(�ㄷ���}�c$���X!%�i��qiCG�񧧱T;iV�uD��޷�]�Mּ;�f���P����x��IF4�F/����؄�n�)�E�X2�$B���#�]�"�Ƚ]��A���P��+&NJ��+�~nQ��%�|4� �� #%�ˢ��q�6����;�[�k�C�Q��Ap#�_B����/n��:�Q�����l5�	P`T�x ����@"�aW�d䈆� ��Y>2��@j�P_*�+J@A�%�_?���6�Zci; �~]��D�����[�Pyy@ B����>Vv�1�S��kNam��|�V�Qs�j.��VC����r�"\;*�JN`*W�oa�
�[ڒ`nC�XI��I����/��@ٷ.���*�ȯ����L��M�1���'=�o�採{��h
��o�%�-Ɩ�x�8�?����y�n)^7y�o��H��Pʬ���o	M��{n���䰪�[΋� �}���(���+6��M��c��S[s4�S�fm��v�E�Q_�?�1\(��AA���-�ߏGU��a)*R���Ľ#��x�ۤ��}�QA����Ҧq��|
���OV��u��6F����7L�����gY�z��'��	gXN���^$]��]yW5bn�[T铍��5���V����H\�Bxe���B�)|:���@=A�EzB����zQ���r0�ݎ��v���1OoU��VaTv9	���q+O��L�v P"�@���k�������N��N����Z0P �����.S'���՘��3��	���7d�h�����fS�'�LJ��r{g�b����&H?���h��&?�b���9�G��z�C�M����S[�a���*gC2M5�J��fM=1������&��	ǒ�MM���+|����*��P��ϰ�f�6�Ͷ��_�mp�v.��:찘�`>T�MA�Ӯ��A<�C�[n�w��r:��������
��ң��&������Oxu��1ʨ#D����i_.M�
�ɒQ�!Y�����i�(�IKz;$��ǝ@(4@���U|b��كdB�`:M@P�eD����Ȧ��s�&��L�o��x���;W���p=b����an�2�RW(�1�}�:,O�q2c�i)o�<�z�'S�SP��]�T���!��3Y���u([�����ܹ:$yܔr�wT�_xO�����~"���X�
a�+9	/a�sͩOlQRL,w��b���QBP�m��Ђ�B%�Vht�&�D"�=���k�fc�tR��6��y��|��q��_E����8���O���fdjN�`�bǉ:���_D�s�il	>5c�FN}���{! �m�T6�$2�A L���`U���NDNB��j�	�Er�q��GV�F�@v��_�9���_��ws���h ١��̾������Dٜӽ�U����"���l�ҳ�T=
^%�|��5���N�@����#4L����!vϲC����˼UG���������L��v6���X�XZT*�Ӣ�#q}�KJP5��^\;��-!�s�ތ�urL*�rh��XL�w�O���J�gxӾ�"n���&���8W�Ж(y�G;��{�v����(�Oظ�/���#"�q����Y�Ԉ�\���"�e�4���x�A��s_��2mu9��;<�����_w�V?�1��Z������ٴm�E�eJ^�?�S�xp9�:$,Auw��X诲Q������<B��a�l�P
������CA_���To��'���v�k
AC6SNd4'�:5`-8QT o&����9����¼jNr�nt�xkJ�8�Q�ࡵ͋��)���[��,3s[�#W�jS��&m"����P����T8,K{�V�fz���6�M��bQ�g˔��O\S�#�A��&��<�����c;qTǪ��P��H�j-��>���z}���s$eZ�J�JF�ؼ�К���g;���P�?;�-~=�w�c�0�+��������ۨ)�ც]�?���?�/��Ĕ�Ey_����²��yc5sa��^�.�g剰"�d���|��dBmG�14��h�A�J��AN3|���#�G��Q��s���:��+�@AvjO4��"��w��3y�PQ��0���*��C
��s��s������'�dU`Kc̫bG��D�=ĆG�^�Ӊծj�O�m���������4p����gnnR4���2��w$��2��C*�=��?�v���,-mą�ĕzh��ؔ��y��mϙ`IH�N��$LU�H�X:+�S�ɳ,��c=؁P�62������DS�����8~�	��:�;&��ːHׯp��T��'g]�RwAp�����R��`zTo����&�+���%�R����\�G�AYL|���]�BWS�gK��?S� w��1��S�3ev���(2xQ��e���q`����N�j�i!����8����<Lxx/�x�R&��8���Ǣ%�g�A.D�x�km��؁y���_�N����4�a�`e�H�I�d��;5�!={����͏��ʃf�im��a���Aɐ(mz�/���nw�S����:Z�	�6~Ef���~�)��(��x��T���t$��I���97#"���L��d�~��<�[��)O�Z�{�+L�e�f���� J��G�<� k·�U�b�A�V��Y,��/4����*�x* �@�$�����0�:"��P_�k��}�VF���K
^aey�7� ��T3`�Z���
3��0\˺AG��W��K�Lɿ@l����c�B{s�!Zc�[��-6��ُ�7�j�GiW�,����Չ�ܯM��۪�m�9{rgs�0���y���X/ |o�f-���2r��c����1�D���nW�[=۬LsFM9�������z}|^[�h!�w[k�qD~P5�`s?M����`Ţa��pa�F�M�Lz��%���$��;�W
Z�Q�Ͻ)=D��n��]�	T�[��O���v��N�/�~�phţp�{e� �LKo�a�}dw��M� Z��(�3 /�c��i]�!��$�5�=�P eF0	�C���N���	(զ���T�|d�̆�gc��]X��:�,��G�I�ؤY�T�$�bm*��R�� �Q���[Sw"ь���f�Z�#)����{�u�y�#��-�N4g��9޻u�?�>C�_�{��B�z"aG����¯q�b��\�ASZ�>/U�1Z��r�h{�Ew�d���K���d9�@�_B<M��7(c�����KfH��?�I*�����!��c.��3��v�%n���[վ�!�3N���$����1��de�f(��6����s����YA�~/��lon�8��\�M̖͒�7��橾H�E~��D�Qc�l�!@��+�'�G���]�e:����U&��T�����LT /!طzZv*7jݷ��h~|�	�'m��I�ʖ����) y�� ��I�^o zN�Vn����M�(Vv�Ч��s"؟��\i��EA�Q�Z����m�N���1ev*U��W�!p6%�|d-�N Ȑ�G�`�6~l��mɁ�BPyCBv�|n)@>����*�8����z��,���JWDp��uլ���������NjӻA�X����$û�Օ��&��d���?Ñl���$���G�d�3ٰ�TգR��z���mD�?��\҇��_g�F0Ћ�o�)���:ȕM��9r��G[��V���L�@ݻpT�|=y�H���UȨ�d?C|Nw�]Av�qX�"�D�z�?ޣ�Q�� :1�Dd2"��;�^Z4�{�IJ����P_�ŵǮ���J�,��z�[��ߝ{e�g��������ko����}w��f�i*�W��.�V!��T��4�?}�L�K9q��	�C��%h�X6]f��R�;`?^!�؂-�g�IE�b=��M�<��(͍��u����h��#n}=�.p�.T4x�ZX�l��Quw����sR�]�[o[���LZ���F��~c>f�@h��n��xI�=��#}5��;"�J��)����6����2x" s�����^4�r�i�����p��LԸ6	������i2ȃ������`�����l��P�'*C��]!'L�&eT}|*���C�ZF`(��;�f��Y��s���S�O����%�
.+c[;��a��w	u�^�m$R�f���B��4�V��臲)�Wʿj�	�t�����]	-��ih��&��4K ���AGM�OI��,�,��?T@��J:���]|9��$.���H�ä*������B%3�a�+U��f-$ӂ����63(ڷ��6��ru%�Z�|iEמ4Gm�g�, 
ϸj~�A��9\�N�p��Y�]�o������N>��o?[�"� ������� �J)�/_�ŝBUQU ���&)q� #�nW���j����w�O~O���E��<=�������xX9�m�M?f_�q��6��2)3y��ͤ^6/_l��0��HvJ`�k��@�3�7lTN��E�}jI\�`J/i���IϏ� ����$o$S�q�s��q3�;Σ?U��1��(S�Z�a[�� x�(��Ke�@f�=����v�5�����ͳI���n��ʽ ��z{���|�@�\;\������솤=ƾ�ϴ�e����w�֦��ڴ-0�ʁTϘ��X���/�uj�t�Y�[�1��#@��F1��b����K��9Xl1?������iZUb���Y@��.�V�������ͅS��2,�����v�Qe��9�Ɉ6��֢7�#�E����r#�;��짛�u����jA�����T�J �d3]|��1Kｽ��Ozma�̝T���F����%�W׃���̞u�[N
ﳠH�J�8 �.�d�V�I9�OGTV��i!�a -��7ߴ�(���[�5��9ep�t�~&��Ι�e��n┶(�l:_ ��g�I���0�䇽�6�z��x��Z@y8ON%�~t�����R6^?v;��/�w
��4XG�c*��+g[bG�D#	���'%ʽ�%�W+|5�6 p�u}��`C�bk߆y�u��L��c�V�{�Τ$Z���?W���{��f����A���n��;d��0ə�Fov(����&:	�R,!*7�&$H��eb�J}�E��&�����5i�����ܫ�d���~x-��:F�іxh-�~����c�ހ�绲
�[�j �C^�a��i"OWݙ��p��hr�nuK�G��E�G�i}�=�k�j�*5A�mx�@آ��y_(�t��NI/ ;�T�Eާ���e��I-{*��<K,�y4b���A��=ͺ�o��鉕��5��m�=���w��(dV�?���h�L�����HG/��n(x0�'`�����%n���Ŭ��q�&�����xf�ِ���j-�ԙi,���YH$�/�PF2�q�&��{��K��Π���R�Y����I�Ѝu+z띅��%�����^�Mc3�es���l�J)�{��5>:o�ojX�W�X
���E(.LO�!�[������f/>��
��V[6�K\c���ai%Z=z��&&�\xD�;M�� s�<|~�]��k�5�x���%�Ij��^!~i����BG�!cn�}yy'i/С�N����� %���X�O���Xd��z��{6�x.�����*kňG�# �!��3��AW9��6:�3 ?$���"�����5�d9�?�&-�U����&4c�z�ɚ�^osmtJjZ�����5!�:��O���($�~	��`�Z�JA{y�4Dh��eSB�B�0��`�O#�A��Ϫb$K��a�����:`�K����?�y�ʪη[���pЖ2�󻱰��M�EK�ݽ3�p���<7���@�S�/�H�m�9��)���G�d��u�'����96� bq��Un:~���ZEI�mWl���$����
��ts�d8-LߊA`x�ygI[����ʤ���v�e�5�B*��S�Y�M��{j�"�2@��!2}l�z:W�.Hi���{=�#<y�����/ruc��S�B���>��P��L���q�f=@�C�V�(��Ȁ�4IÄjL�(���2q���~jv�QBQ�Rj<���ɲ�L�t>��޿8���_G
��\!�1�?�[t�O�#p����5T����ˆf8��=� �E����#��~�1��@��?�
��z?p����f]Vu����3�B3���x����<��U��yZb$��v�݃���D܏�Ѳ�O佋	��8f���&~̲J�)��o�6>0���[.ӓhm����'-)�JyC�@��C�݋n�X~���&�5֎ɼ��.�V�'+���9��D���@X��(g�H��g�.##^�E�}�Ϫ�3޹H�U��M���(Q*�ڃ�Bm$����9��4��/��y�!���o�?yH�Q���6�i@�'�{0����|���R3����б	%��ٝ�Š	*�L�3�/v
Ye�nտ�V�Tz�}i-E���M�)��h����Q��jjf��ʜ3���<đ�u�	��&HǱh�F3�����g��.՜��<��`�V����C�RԝM���d�=6�CM Y@UYF�f��u"C����\�T۲�z��~&�)`}i�v@�g6aJ�O�P*��~OT ����Ç��b�y
���e�(��P����u�⥞�g��������E�AN�%e&�B��>��|�g���c�
���%�E2�B<؇M��\a,�6�u-��s��kiu��tU׃������5#��b��J��
����H�ъLb~��Bz��B�	�wob�Ժ,,N����R���� ��c�~��F>@K2���~7:��?(�� ~��j:���Ůb�������sV�G�I�rû����ƁJ׭F�p�n��qQy_�ى{���v?��D���3�X��_�y ������e�!�F8)3�u�_7U��z@��$�5�v���=��&�J"��bVupY��R㈏ɑH�]z5:-���j��̅��eBs�a�nN�����I�p�Ϟ*�#����Yh�P^5���R���q��/ր��6���^"�pzIH��Y�`4SA-���� ��J�k���+�i�7�h����F8�}���[�!�;��b���+�O`�#�#0�-!�#0-� xd�u;1�iS�ֲ�"]� j;g��H�+�tb���;���)��/FZ0{���D	���ͫ������-��u�m)�擒���?�H�&yK��9��شwGY�n8��&Z&�Ĉ��3,�x=��s��S����|w�wuH$r�>�s���H*H�0�:�A����4�ix���=����{�Mn+�W�:5L���B�ov��"�&�r�o��x]$_Q�Mҫ5Ns�f!�?:�#��#T�[�G�����翥+i1��+1�"�����;K��e�X�E]q�w������vû�2�7�ky����S�j[�,�
���y�}���!�Lxi�G/jj�?z"Wa�I��i᝗Ei�|��OCq�aݖ!�E��Fo|�,��V7������+���3�b]]s^��;T���P���8Д��#�S ��I������ ���p�6��l�Q/���l.��mE�2�x<O���R%�Z�����{C�]�a1p�<7�R��a2��&�{[���rަ��@
�I��u����W]�E+��~Q]ʅ�Ĩ��׼XCj����A�yC�Au�������rz���n����%�
�����r�kI�>�c�Ù��Ga��F�Y�Ol&��)�X�H�wV4��%R�6�
M�h�ؚ��)����_��ڃ�8x����횢%�f)=�na��_�"+O@OF�%6"��#�C��vs\���h���k��Hn�X+��p��� ��#��ZE�_���͊��a��^EW8��&rQ˞�&N�gu�מ�XnD�� �S��pD����� @�xn�f����q�x��O�`ɣ���{�e��=�ʟ�NqI�u;���c�M��5� Y`y`CG�[]p�BV䈕��9���,E����ʿ֦P
N��y���"�"��?��P|O�f�忯Oc���ae�y�P�If�2h�3'����?7�E�%��_`����t���|�5(�	�o���%\}!���Y��S6dM��_8I�[���wM������B���W�I�lŞ��S�����ϰc�SKs8/��]N\CȆ��8HmRp�*�)�]�����%�����w� �{�ڳK�rz��%����(������@kڏi�ޛlo��0
J>/�c�<T,6�b\Oi4Q�4o{#����JV��ǍM=�X�\v�������y귧:z�2gS��Ě�)$�y��J���$���q?��q��~AĴ�$R�Xe�}:��z�F"�Sjҫ����hm�_�va(+s�s����:�|���NN��x/�j���'�c��+N}W�է�me�#�TG��2/���)ܫ�d���mrI	����F'��t,h�d�2�ń�-�DBӂ�-��7�샩�Jr��`:qx9��s�Q�޽ඁZ�k���7z�b�g�y4<��M7�?p���� p&�߁M��r���8�`G��y޻
��9���������l%'"q%�f�{#��OQ��,�U�h������R2�D�~�C��E��vYw^�Y49�i�sR���Y��m|`j�׎�Y�<���>��5ZL���$ӆ �ɣ��d�����M�������0��&e��QP4�{��Ѧ�"�Q��7>mm����8�߸#�8Z�#gr��Rzo��1��}���)��Ro%�TJ���e�@fe[�6�P'j3��~�fN�Cιi���1�}	$�Aq�����O�� ^6��J�XbȈ�g�x�au���|��qVd� 睝W̃S7���7G`u����1����*��o��L
"�&uK5�r�Z=��G��J� Iq_Ϲ��d����2B�
�ZX�7�p�.��n�L�Άxvd�a�p�툚j� l����"��%Q���\��A��`��ytD�N)A к�TXd$N&Љ���{��t�K�����/G-��n5�,x��.��2a��0y�?!`p��~�PY�{Txf��0L�'6+�W_[F@45� �;�}Xi<��C�'�E�a���o
�Z������?��%ŦY��-�k����(w�����L|E-ML��#f}?��6��'��I�`����(7Ý���C��0?�&�}7�? Z@@�;��f1S�A��X�1u�c	g6��LR�����H���!��r���fR�Bf;2i�K��ex����(V��d���ϳ!ku���U��-��
r5lb�rS2	�͖�A��u���雜,��K9��Ui�H�eLKqO{���`�������#�M����m
�J�����#}�5��������X��I[	��9 p�)��*�4��� >�.s��}-��$mC}���>���s�*:��!�&��o���~6�6-�AX�J�������і��]�N����,Iݒ&���
&�XQ-��9!lBk�x<���-�ɡ֊�2p[���]���<����|Y#�&��Y6/���~a'��W@�/�fP~Nc���P�����"TD�gD��F�[�"pj=��W����6�����\���u�x���SHU3w�(�M@ì|�ɯ�N�9C�[�X����<\��O0ۙ�y�}k�ƪuh������4��!��:���>Xֽ�99���ٱ�-�*�I��1բ����.�R�`�ݱ�*��{��V�\�[�`����oQ���2��Z	�:��^��&za�^Bŉ/�t-�����������	�X7e>��#Ub��.��:�_C�g��N�cIfk&d׃��]Rk�o)+��Aoݐ�E��f̹���[�r
�;�oh�������d��"�S+c	�c/��i_�ߖOV(T�!D�����(F��t����p>���$ˌ��נ@`��6���13�>�4ԫS��:�[Kt�W�����8Y�Չ��"_�;��E�B&���*�c�n6��*ȾB��M�Sl�|����� �D�=�byŻ߷ �ݗw]R,��I��ʖV% '/K���L��l�K_�a�	�};��`����L�"?�q7��S�c�� 
2��,~�뚺�z�ٞXg���[�����g���
��!�mz��h[}}]��J���12iy�z1�gj ��j���-h�Qw�3Vu�ڂ�V��m�7��Ճ��<H�=w�6nY�a�����Щ��aY���-��j���~q9y�OH�y3%��&�+�r�}�늉% _�2�P��]su��)x��_����\�D�-�̪7��l~�$�R+� pDT���v�����T-	2�?�ﵖ��i�f��b�������Ug��U���Ӽ#���4�e��$Ѡ�V�ki+q�l�L�A���#l}�?гMЉwK 0��`��n����@v��1!�;��ǳ���f<�)*����mQ��J�A����
�8k��n+��̛�����O�o65��A�C5@�m��AWv2�Q|a�O���X����-c���*��w M?Ȩ.�p�.�K�e������������@�#w�a�����ACQN��������[ 5/e���ɑ�+��o����CS�N˅T�,V{A?c�@ܩP�	P�j#	Σ��F3��'�&�&E�B�������Ddd�eq�paFۀ�⫭E��WO
�)Y�Y�8I�8,��o����AB{wk�^�w�a��P`3�Jѣ�%���E�K�"�a�-��e������@+]!��rn�����f���p�+��!h�c[6�?I��]�A��?� ���4$&�B�f]�pC�b5����e��l��	B�t^�����Mޜ�.�zL{��e�f�9Cp��J��d��s+��a ����ʣ����Z�+o@�J�+���Qf�D_��Sݼ�P�<kdC�)81̗s�WK�
@5;����**$������5�Nmyu���k=l�%�!ma�.�1Wn��.qX��S$H���^[CN��L��̱f���M'{��ϓ��g��Gف}�=�p�����#},D/�^|#��Z5m��C��۸5�xj����" s��7��� �a���n�c�� �iL��Q�^�Ǌ f����:�!j%-����q�3�c�����A��i�ʷF���@�~Gc �42��腳�'� ƈ3Gӄ��.R��^�Ҩ{@��e�F}�k�9|��qn#����H�P�V3r�s�-nZlj��Ւg&?j���B��a��;�W{0�s����Ji�Y��i줾#6E�C�yě�����Ҵ�?2_���'ݠ.�������{@�T��C�TB]�&�a֑�J�A��c�`��`k�S������C^�Rx��]w�9���� I���͉$�Z�\Rc׊�_5	�[�߼�:��*��P���\^���Ze��}�:Sb�D��s'j)�q^��r%�^)���h�G�BR%.8���x%�Yl6��;�L��)���j�@�d]Zk�Kb=9�.�o���><�7l��r�W�#Ic"�؁[�R������Kx0� ��)�x~���������7�~�(BB)�#��p_G�<��0+ːė?d㞘�Dzs��}��.e��d�q��|�5 �e���K�3m��p��~�N�$�u�����'WL}�Ȁ����){'��ȗ�2�[Q���i�h�ᆮ	7p1̈Y[�D���܊=��.��a�ݸ��bYM���}�^c���CG`/
�~'���Q��=�����Ij����%�6����#��&�$�Ҿ� �1Z���!��E���S��2��G-~*����C���Z��P�8�,�h�:(�3 �F�øD_�S�	�&-i�Z��&Uy�/�W[�t^@�Q<ɬ>S�zy�@˧,8@Z���ݟx�d��I=���u�N���V}��kXa�	�Q]Du�E�1�ktw��h�O-U^�3Ǫv-��j�韷Y^�>�M���+�q7?���:`�8�«��O�����E�gd���k��%HPo�,�'%���7Ӏ��AM�s�ʈ/��qbRCN��b�K	z��� �#��� ��M��#��ad����l�2hCdT��]E�I~��A2_�z�ڧ
8or��8��*���������[�b�:ej:��v�4����>���v��z�;x�O�2ͽ�Q�UxyV�:;��8�]="!:�
p3��RnS�}����eY`0-l��0�+� �?��~8�m��|[XP`郯�O��7��k�,/�`]�������������W�A~	@T]{���*��s��W�<�b1h�����#ɰk���-���ܱJ��Z�s!��5i�S�w1�����@Rd�r�X_Ӑ��<~zS��� ^S:��ʍ������
��2��4�&���j����R;kt�y�H���?���a6B.V%G��j�C��"�E���:?R~%�s*p���"�����N��Hq��z��w�I:�Z2}��VM8J���[5��Φ�� ��F���ӈ��\�d!�h�F��%y,	�vWq�	 �]s!� ݏ�F��]��r@.�6��L2��p?꭮-�ʸ6�kUq����a�@V�F�
ԛ�Q����1���ϝ�����'��Gn�@&�q����r����wXU�0)Ϩ��Z�~��Y��M�f=D=���� �@#@��d�	�_䦞�I���t�Tu���g�Ep��S�(�4u�=�~�ح�ݞ
,d�ʳ�%�Ҍ��$�>:��W�"�\X��f]0m�j�D���7պ���C��.[�8%h�Λ=r�PfȪ�v��R�j����g��r:��AD��ć�brP���h3�j�k|����vU����45TJ-���(�3|����=�iE�]4��6�$�tZ.�ћ�/4�vȨ��p_�blqސ:�|d�t o���^����k�H9%
�h.$�n,CҞ��dD}X��>�$�[C8>���X6,���lJ�K���7�>Ζ����;C*�>\%R?������̞1� g��̥�����{!��Y�O·����� a��)P2 �AS� �(��u�^�ʜ�#>?B&J�v�զ��<\���1t���"����6�����m�m�� ��%�����ڭ�ӂ�9��I��P�L�:�H��3��R��=s	��k�|?��v�;��M�<��I�� �,�1;��9L���^�\&��B$��ԍ�|�դ��I\Z�`C�B�2 L#�5l��*��ҹ�� jI�"-do'�V�Ⱥ�ջ��#QN��
���k�]�q��/�{������
���,��9�/4�jm(bJGI�濥db�0�	O���L�W6&Ni�j2X˅ǳ4��g^�A�7�M �$��F���9�3�����\O�_�����d�Vy�Pt�L���h,�bE����n�ol#��.m�Ce� ��K/�1���c�F������ś��y΅ܴ�+�c=[畅�B��OJ}���ٔ�Y#�&7�l�1�[EC�.U,?[H�x����]���12hU�Mh�y�����0��j�U/֙���^�d��`0�|P��H�#[�>��u��Qe���P�ޮ��<������}:ц[���
Y���\���>?X�f9�	"��w��\�.B�����9���������h����[�Ƣ��@�o8�i֠ӏ������ǕK��A}��M�����%�����0�Q�F�\kX��N��5��*�=��>��ww�xx��A�Cu�(.[ɣ�X��n���cF��ס��[���f����"��jy�>h]~�C�pG�tAU��lX�j��}RD�k��ܨ�iFˍ,FB+%iL_�ó8 Eg��W~�i1{2O�}W*�����Z�6���k8��L��L�Ľ��`^��b���-g0)$TвA�)���KO}�]'l��lQ����4H5��_7L�ZI6���Gd���q�Vr�yRj�$������F�;���!"�� iòӓ�A�{���� F���wr'(�dwOxg�����af�0N{҈c
)uұ]B5jy�0B�KJƯ7��}�P��T�t�dF�\ޣ�G��%1mD��[G�s*5���L����v��h�
L	5Y~�zц���g,P7�H)��;�X J;R"u��>6�;~�Rdb�j�}a}�[�w?KZ�4�+�-0�&?��:�I��ri��<�4�R��ּ����wW�^�����J4>�&������e����qA����e�V���Z9wVs!8���C�`�����Z�83��ߵk�B0 �(������V3������\��N�� Q;/9�`p��TJ~o�H��|���r��eI�FDH��Iq�8�r�Xf�h������
���LkL}.d��wi��ޏP��W�S�$|m"[X �a1|�*X	anh�* n��F;�>�)���ʖ������������Ӵ��^�.��QO-��S�Х	�q��AR�Y�+��4�x����(�/j)R�S��ہ �M؜M�H|�	wj���!X쥬�m۴��q�Զ��f;B�"�.[��{�P�����`d�I����־�������-�$t^Q�!^2-���͝3b�^6�z��X�%<L�z3�o�!�_� �
�0
M����Y�
����0��_�
��vH�'���ASz�]��3i�ns�?��i4א{�t����]�����Z��cs(�I��<��W�N*� P�l��/M�ީ�r:/�e5�J"��|�d�և��P}GFN�O�� �����|��������(�؝L�#b�#xs���u�
�<�Ź^_ȜX'���<��N�����0��_P�.�9[��z���ݪ����(�1�����Sh��"�/6�J����Ŏs�ת�_-�^�]�����}U����?9��[ M�v!-�Q��'����g�W�U�I���
c��Bό��l���_eg��q�~��l<}�"�o����Ytb���b1"p,�b4S��\[w�
_�3��Q���U���;�|�Y�D��ؾ���E�<�/kH�x�X����Yi7���9��?��@L�����m��]�_��l΁QHo�53+��qR�>	��˔^�2�����f�d7�َG�I�g�:�j@��}#�
t�j�y��y�;�$.yN�8IlC#��)�s @C�T:���-���>ҏ���@VW��=�;4)Y~��qr"&m���oK[�Mj��4\�$�I�����{�ڧ��Rّ�a����!��G˙��>y�4N5\��y6-���\�7*��L���CU�b�_\��`���5�{|t7�^fK%��>{�.��\g�3�穃	~�V��өXșy�����y��2�{Ğm�`�����V���A		�o���<��Kb�JR��_i�5!g�?�	�Nr-�pQ9м<��!� )n�z��'Q{�?K^@��B�����&��0�d��% g�c�0$	!(yE�w=K�����8�|_�ʳϨ��1%m� ��-b��9�fk��ᩯpY�����`�ue"�>�|�k}�}�~�����/���k�Ba$׍���֛���YN�Fw��MF�:v�&Տ�;ɀ���V����m��̜�'>��W���i��B6�t�2L�1t��4��x�A8�c��ɏ��u�����Ȃ�*�6F0� ������
�J�B���͗nM��*��h,�?hqGɶeB��u���E�c����-n�h?oV4
�"�����Njɟ��n5�@\�.�I�h�=�����Es�/`��nlK�;X<�A�}3����Uc "�L@��D���{�����齵+�rf%t�(Ӡ	W�.+�*���@�>)�`9�B���ƍZ��&�-�l�?�_7ɏ���fI3�M���!\�ֿq^�O�D�L�z�ς�z�OBtQM�J7���:;��>�����du,�rc��Sf�Ax�y����
�F�Dq��� �pC� �����9��4��h/8�j\@D�i�'�z��Y%'X��^[8
�����[ē�9�;�s��?�&M�В�jS:C]Ѵ+��UDPB��L�3��b9$x�{l��p��=V�&��"���j/���gQ�DU�}J��h5p��L'�w��݁7z}ms}�Y����hj��L D�����D��U��5���sf�ҮjP���)���=��؏��7,$�"ޫtz;s�ʽ�p�9h�{��gG�*�F>��2�$�^A��%t��T$|%�L.&��\�w^�x}
�$X��ꁄl�����ƚ��X�1,�#!S��ž{_�ƃ&�؄��in`��/oLd�,[�GEY�q�a4T�4N�Y�GQ��c�,;ձ�h$T�m�4��JQ�e9��7RZjx�7��[Hg�i���G���ޖ��c�� �b�<��毧Cm�1�~r ��K�qs�3�`�d�1e-"��u��
GZ:tym;Oq�>���7�l��3B�$<�4�L�����l�Đ0�"�+�C�@�7M���sQW�}5$o��䲷��x/M�֥�c
����n�gE���BroS�oc��8 k���z����I�>�.?��ݷh[�����L������k�Z��WcKnm0u9ڀ͐���+�&�0��Qbwi���x���OY�٠F��x.�P�Mu��U@�>�F;g 5�x���=��&���
�b@l��q���ޙ��3�Տ2�H�r�(�u
�D4؟S�zpޫ�2?X�b�ٹ�퉗j��4ܛ�	[��+�p��~U�:s��$�K�"��|,1J�ؓ�-WW7M�W��֌C�uT�]S�z�L5�,#�[�-5ޖ���v���Ӑ�W��l�fe��2�!4dI@��H��w�ȳ�uv��q���a8<��IiW?ɼ4�t��?�w�$�Ķ{�����c�i��b`�L���,fI����rA !^ 5�%��>բ��+��?bF��$�'����� Q`O��'0T����[XA\���pP��z4I�@�m��?e[���\I.��c�)�q��I��čɁ�@A��)��/�*�4]u��͔��/�דak�u�t�bx(�	ݏ�x��"�E�e���%���{g�Z0̀��8+h�c3��fE�}MUN��{��-��(l�e
z��ŕJ��:��]��Zl-�f�]H��Y�h0ld����xZL�Q�nq�!�#��b�~��%@�k���w���,�O���]���
�7�}+��.y���4JU!�۩`� �:e�Ҩ�׾�,Ai��$w��@�^��-��NϬ��j\nQк�����N%��W�\����G1�7q�`G�+`ڭn[Q��qza=�k{~jx��|��*q��~��7vw��Ԍk����:N2w�^V*��HӤzW��;�ݳ�<����aο�Mդ�iij����ٚ���gʅ�^��	����P������@��U�����c"W�A�sѶ�nYs�=�3��.1sP���8�9���'Ő�����a�!��Mi(_�9�zp/�V�]AU�v"��b޹:A��l��l����%�ȣ֒E,7D;��FP�]]�I����E����>ջ�{�o��vl���ٱZ�J�]k���1�*�	���h ����͈u��bŰw�^].H������Q�$'�q�l@b�|l���~�s|�ԳY5��i����ޫ���C���2�+���Zu��C��D���?W/��Nh��ź��Q��>�C���A���BoҰ֨��Лܵ��E'��:S���bF*����I��,n�
*����q����TRb�i��Q:ˀ�qfSN^j��pf�L��t��W�]�U>�pYG��������K�ZU�4�
���;�\s ���`Tu��Vx>XO{�O%˕؄ܐ��>�¸��<*4�,�`ѭU_��"v7D�§�Ir/�f�����GM���tu�e�%�N�wFF�x,/@N��5�y��fn=�����8ʗvQ�5D��t	9	��33�]xj�����h@����]Ц�lU�
�I@t8���9oF窘�ko��b�����s͂E���n�4���6����qޭ�`��}f��o��X2���`�h���T�ӷ��"����{}����v����0��9:[U)*ot���e��QU�.X���g�|	�	����n&��.���`G���S��\,^�O��4<���Z�66"����������-b��Yɇ��"�$�w�Ve9������"�r��U̓��P�Ǹ���N7esN���ȹ�QN�����z�<���}���Ā����������T|��>B3O�9� |O2a��A�I��jߕ������Y����]���SM7�j���bǲRר�̷�$�7�:77I��?�}2ߪ�Q����:M��*������Hү���} !.y�
�kDFF��"hj]Sj\L}�~�6t���3(l���kf��G8��f�[�+H��RՓ�7=M�Z�7�C��uo�N���fGEb��N������~@=�Lx6�}��t>��0�.	K��\lS�"
%�W�
����C���3`̀J`��	�����W��U�vاJi�rRi�c<xn�<|y1ЧTAJ'�t�"2{��(�?�37|��S'蟜iH_uS�3�����X�I�޹�ޜ�e��(���#�\��Uwi��(;P1âS��tYo�І_ø�{��aju����4xK��^Y��HP�I�U&ry�|j�?��C �QXuB։��H������c�;@-{F+�'��c$��� �c�6&�����GT��:+OD�����h�B	��j�qҰ�]*��Z������}*������������3�:�~�@uj�X�p5���В�#k&۹X23� �^L4擂�>`	�S�Ή<A��č#hP \ʽ�2��S4l�E	�t|8�^ҿ��ۊ	1(dB��W����IO�du�B<�C6
�?E)|CԞ��nRD��z�5.�-�`xu�x���"��3��:_��)�`�O�N�_
�W�t�ö�*0��zM�T����IU�NwD��4���ʝG��gMS�1�*�������#�ô;0؞ϑ�ާVц�<��5�����I���`\�|΄}-�@X�C�_�@��2�('3�!��Q]������>�D�x���F.�%��kW�2WB����X%C�l����}2$o�A�=lX�a�����b��Ż0��k9�Z���,��(�/�6�I:�T����t<�'��U�=��j
���0[	��4B����T���J.Ȁ
9�d]<X����\ر'k�K����XX�R�S������BV\܀�t�csǄ����N�f|�g��:W�(NK�IPy을��b(#�n�y�]��v��꫟�����]&q�d�\�{"OS�z|�ZG�P�'�á��n����w`�����y�i��k^a��I�����T\����l?�����h�u��X �����X���қ/+�!ȈW�7�c�:�2�ң�6����М�m,�@d^S��F;y���)�t�?�ѯ' c��Wq�$���3�F=b�[��t�#����4o��0u$�m��1/�:��]Ƅ����n�6we���,�<\�c�];z4L���i��d���4ڈ1�o�p���^�pS��v���kNI7h�
IH���Uc�˚[:����`_c(M4p$d���|1TҜ}u��(�N�2�ڂ��^��e��H�0$y{ʍ�^��^O�m8��9�����e��46����l����*�d���=A��):�pc?������OE~5���W<fgP����u�*�#M��v��tP!�U�{�ü���?�p����c�E��s�+���}]�J������MMm�+~G�uHB2���z1}7�8�=K:�U%�Q�}5���\�& ��h�
�
:G�䤍�O&�ؖLօ�@8��eN�9��������P\'�sGIRM�kH�����$�f�~^��ʿZ|�9�ʸ�0�����}�R�N�)�"�rǯ��$L]͂�Sub�|b�B��"�_��*!�j���J��x�[�&����ĉ��^���rS�O'|d�ɺϘnQ[��7�B�_��ɸ��lHX�E�}_=��)���a��j�"}��m�*�+�J���v���*�D�u΀~��-��� ����,Z^�V��gYn�/u3)t�!�C�����c�7'��TP�(�YrN �}�$�k.��v0b�	c�E/6�G=3W	��#c��Y���æC��%B�B8r>���h���o�Vqd�ڟ�q����o��c��>�Ŋ7���ݩ���Ϥ�Ӈ�t�S���:�}���%R��鼌�G�A��,gF��	u!w�c���Â�1#@�Ծ���������R�>�W�3vQ��*��$٪� �*.�{E��G���v4x*��m����ǈf�7g���#m�8���r��G0^g+^A}a#Y^�:�{)��ī8N4���wi�L���0�v�<��uP�����>=�W.����/z�.��?�IF㏬���I����>W�;��R� i�ۺ�@��8�V9�jz#��F�W��;Q@P�X��!7��7���z�0��I���A���Ɏ��d}o�N"u�~�\T���g?�����:ud�BJǊ��A��{	9<�H��$P:��R?r8������'�qmׁ�-PB����r������Έ�񿶤�#uh���̷ �xךZ�k^��m]���[~6�i�+G�g�TS�!�`R��Ֆ ���sZ┈1��ҳk�%��I�i���£eN�zW���R1��b ��o�ߔb�Y�5������ɇ�Y���%a�Eޙ�W��K
<�{�lz���D\Ի��U�MF���]T���r�I�2#�o�������W�]�:wb��YN�c�6`�5ƚZ�i���槑�Mk4k�����K|�M[�L�>Ba��C��@��q];2�ݕ �5K-��)��8���p�멑9��������|�U�=����ٷ�����V��A&�ǹD���XW��_��`z��f9�4	S@g]w����1r����ˎ��n���"?q�a�Ҍ�� ��P ��w�t���(W
!�Q�����7�*ɋⷘ\�E]�0�&r��x�q�,
��E\f�N��hd�JP�RL�ëhΤ��E�#�H��`�s����3b���e[��@2%������oz%D̙̕���_[�Қ�|�l��f�DШZ�I�A��z�/Ym"C'��������ݷ/~o%vs�S3};J��:Tџ�D"nFs4
��E�)�i��J��Ùe:Puלz6�dc�mM�;xM��XOAf�+=��()���
k�nQ~Q)��(p�b�@Ɔ��.­��oB��8Ǟ���ҽ�b'�O�7�ؒ
y��m������M˓�vF�m�=��C��HZ�@���4(� ��ȵȚ.��dm��<צ%Z'H5@e����e� N���Qq����m�,����o�' �1��Ad*|��O�:�?�k�j}6�o��9^������u��Nh\�?I���T8,{u���Q���Ft]��i:NKH)��
��3;� �OJ���K�@�|Ђ�΅��d4rhذ����k�3����w�Y�"�ME>��^�ff�˖�E,��������u @�����w$�w�#�u3�9Bƫ���]�˞"��=��}��L�(R��!� 4�һ�I���$�1_���f2*	F�ō�^c�8�%· ?��Q���Ҁ�>��̓{G-\?�F8e�䠳��w��+/��*<6�ދ/�� ��m��Ƞ��U.�R�l���a꼘�+���/����R �RK��m��tk����do�F�8�\i���Ȗ<0s	���3�0�%=�[n�s\�?�1L2�X:�Բ>��ꬢ+�\�Y�t�gK$�z�DuXx�b�͐�֙������|J�G���	�V��=Q^��e�.H�㠗�;���XJ�/&7�.�� ]X�sF������*ɴQ��m����3�7t��믞��[�BH@���U2��F쯿�1�@_�j,��ӫ�'��}�g��m���~�����Q㨘� =�?�ݨ[�"v<7��rK����"A�df;S�U)��^�d��i�<�!����0/���S8@�?�Q��84U�Lչ"h��W��U&�C��G2��rgXi�X��^B�c�}g���LQ��kHT�L����T!K�,��l�)X{��*<; 5]�!�1�Ȧ�U�����\���.� �Cѐ��3{M?)�R dD ���V����5/�"<f�5���r'��C���u	�SO� �x�RO0��&���Q��Ay��KFq�?������=���o�r����\��6�c�XHm��PL�1N�J5=��L���V	�hhY��L2�.f�+N7i��*���D;x]���p�jz*�8H��]�����\b����@��#t�r��(Z�
MH�@��Lj�z'*�+�Ε�T9�VVt�/�pX�{#�.���`f~o<��F ����𘕳vW���\�f_�d'.��8��3fF`P�o����v��Ka�p��)1F�|謑�[ai�F��@��At>P���O���^M�e�T���ܐ9�G=�󆻈�18¬^��p߆���Xj��B��j�5M�U��v����^}�����m��������6|B�iNDv��g1ξ6�/}*�����[P>P����ڳ��QlZ��I��U4Hǧ�Se��9������s		<���S� .n�Is-�aW���m�']��z�&�U�<%WB"�[�it�*�-����Ȍ���U/�τ�T�e�<�WؿYZ�׭:"��!9�,ko��=�%P���Go�GR�$*���b���}r�rR:5=,X�}���'H杍����0�����T�iԴ!�@b�z��[*��d���&��8:�u�n��U�&]-�vO�#����ڟ�Zm}!�A �FI��v��x7�.=��Ă�x$-h���'�R�����.��u���~pt�I�8u�����Ш�9˚��|���Ԙ���^:�Zݏz�n�Ɍ�o���ig���W\���7�$�L��Mxtb�Wk�?�O����&;vw9W1y���B9��b֬��[ P�����U��Pk����4��1�(As+]��̿��0^�=��R�Ȏ�q�*�p(Q+K����.Ƨi�"�N���>�
]�#�_Z*A����
z;c����_�%l��t6]���H!oּ�_������,�a1���,:�ʋ�c�Q��b7���쵢�5yį<��L��tVy�f��7���1�N$�����o��ҝ����8�+/�e8*-mo%��3���%�n�ٵK�jieM܇�A�����Y&=�	�N�^F&�ΔGq�.=��G������\y��(�tx7�.�:�
87�5+Z�4W���x���/��m�<��a��z�o��5�Ĕ��EyK��4��M�-΀�ydkc^�����7L!�"�3�����$~e۪y�I+�g��d`�ڲ����x����~���/�*�e`��7D��Bè��|�^���m���Y7�U�u�Xs�t�RS���m���G��#+Q�)���]��i�ũ��Zk���s�Z��L�'�t!�ʁpd�&f����Mi�BI��@|�i7�`N�^�1px�����/��-���3|f�*�C�<����&�p���Lf��fgl-yA�״"t�Ò���I�w���Cb�v ˜��G��D��#i����(�����;*#~�4��`AdV��x�pf~��vx�Z/�4��S�o �D)�џ�[�V�0Ė�,�.g ����Nv
 ��2mo�<��ޡ�}n�ł:�On��ri������$��Ab�/ΙB�*��ܨo����u�l�K���������wH�%Y���.K\g�*�!F�
_=�b�ڠ�7'�u�
�|/�A�h�9ߔ��ך�ea?A�x����`b.O��CU�Ƚ�7ܕ��u��Ytʕ�b��)�4���c�A��q��i���Ab�"����������yXI�,�C�<+n�4\��g����'��j���<�W��nէz4�2���FY�l����yi��8YU��DIh�Q�q��ɭ�]�y���0a5TX�S������#阮4ߑ5p�#��g��
 ������ /Ѧr��c��~W��r� `Uy~y�(��kM�ݛ6I1x�։A5/����.ǈ��'��ٖ����%i�0�/6~|F�k��#�E��j����W�{�b�!�-����@z�,/��y�Q����isky����=�@TE��=�B(�[|v�'l���G�B850�-������XiY3�G���eb���4<��P)ޠo h�W���<�}7�m�m�5/aӌY	~��͊��ͷˊQ��W2���c�gU��(T�����Nu1we
�iY\��D�@a)���� �����̪k4��i�ɒ'�I�d��+0����ZN0�g~F���a����Q9����d��i�3u���Sj �U$�&�i#fd4^c{��Zf*j"����9�d����L����2��{�C�4�	�#��O��o$Ƅ☿��>�����,�*��^G�l3�������p���L#�?ɩ�j�z���S|�ۄ���S=yc�+����
*��ǩ����V��_�G �R�7觷�0�uq~S'R�<Mh�0�M�|��ȱD<�@���f�t�
��/�~&?��D+|��a�_�uYnٵj���޻?>^�M5�oQ�dΑ�#�j%��!k�A�����P��k�u����.Ȭ~�=�!���Ѿn���{����T�B���K�)�����HtO9p��r��(p�3+��8~rO��q#�9AwG�z�6��� ,\���,�vY��drfv�}(՝��7~�`)
�ֽ��[q� � 9(��N�<'*�uv�?w[r��~��l{��䔞�l.����>"�4�-�Q��~��x�ʎ�CL�i֩ąd'r�)㭤V��'=7�v[�4���8���-<�	����Pb��|KV��"tO؉d�U������DFƘP�]���Q��̏j�
O�4|U�7柰�}�"x���[�E��|����/}���:2)�q�U50j`8\1���,*[�`u�V�Bh�ZXb��"�rs)}���>�]{= ��L�h��G���Yep=��=�>�H�3���Z�n�Mэ)V���Y�H�N�X�i � �P&������x�W��*��a�c躞�4��m�*V��R�|�d���EI�u�_$wAO@��H��*�+9��LG5A���ؾ�na(�����R�H�H�qAb[q��J�Hk� E��@�77�-�><���}���!9,��#�AÏ��ј%k,��c��
��~g5��&� c�������jY����Pi�I��e�`�����)����ϘR�\�f��bK�K���<��]�(�K��UܲP7���~-]�_�	)������SCjk���9y!�x��m>]K�^��D����&)^�v2z���7��H�	���:��*�]}W�� Q�Q;����h6���G[��~�g*y`�;�m�����D�]���g�ײ���r�[�a�O���|��c��zTY/��M�!�KC��[�e���Ԙw=��6�1�5q�/�Ym#��М_�r��?)��j60Vg���7�I�8
4/��z�iE�T�ˊ�����X�e5vt�Q�巏P��nK:�S��"�\�ս�3�{��G�`{X�mc|�M9݅����I���]O���K��U�)�כr�*���.�D�+u0�K�=r������ĝ<�@a�) �R����T��9�����:n�N97���{��HR����hdbwZ,?�M�b�L�г������H��F�OĘ�D�<^�<ȱ��{��/9�G7%�i�����^�/�O�Q��#sK-�@f7�!D)Ɯ�ߦ#@,Ӕw9+�J&�l�ǍlRw� V�����I���37`�W��~�b&R�����/��b7:p]���I�;H_I:d ���0�n�h�ލI�{��x6�Xt����JU5n�yϟ_٬2*9{�<z�����W>�pz`�5�N�/��.Fv���4vT/�R`����mR+@���Eg��5xj6o����1[���+���*�Quƨ�s�+Qm�Y@"$���M�Ӫ��'C���a;_�I�	$sm�~��/�!~���^P���	���+�:J��W��]�%{�u)��d���)��Аʿ��F+4bI��^�Y��0�<OҚ�tb�*�ukem�t� mX��\j���EԒ)�(ȸ��M2n~~�����uU���g�Nߩou�In
DΪ'j�#PQ�H�(�eh<����$�|��b�'ή�D�wYm��|ܻ�H�����L�Y� �{��?s�W�*�eޙ��\���^ �a.5�q�{���u�z2�sf�
��v��͝� �D(�ft]���@��A��q���RF�>���;�>Wٻ���E���W��?±���S&�: 8v@r2�y&�T$;�����*K��Њ ��O����1gC'g��d���/z����W�:$�0����=��%�w��hG��$4�oWPI,2�	��̹t)�ۡ)�8�4�����k��~v �
�R��,��<з����>��;�ϯN�����T���X�0��$Qo��ǹ+ׅ���"�}
��h�!�����X�{���i�}�6s|c:�q���A�Z:�`�PmD��ė *�"5i��v� �
[��F�q�v�rT�N;�-.�%̷Ѿ�1�����	��%q�ڏ��J�v��D%��a��oD\��?,�]��F�sA�5�e.�"�rt�t67��,�9�o���#�xVa9��)W{�O,.P(v�]O{/n��ɳ���Ȏ������(����l�]v�����u�RYK���ZI�r�ޠW(X0=���$P�6)J���o�q��r7ޠH GE���Hl��#�f��0���6�ߞ�>~~MF��N�e5����&���6�=�7�٪�YT�z�����I_�g��<j~j|�t�2ػ�W�����#T0@cv��Ef*���p}O�bR��4��-��h��-��<�X1��ze�R�ec�� ꇢb>U)���?����4,�����~���߷+�아����#���b{�L�: �`T�܁�bX%�^�UR9�,OTOD��#4�O���&�+(�z��Y����y�K�<�[�6�)��XA�$�`40U]��C�F�ç�G�
��-��I�.�g/pvr1�t`�έn�Ԟ ��V���{ḯ~�T�l�<CJr\|�B__MbU�30��F���ߛ˓��"
9B�2���Ӡ�Z
�yd;��H�9*��N	�+:}T�!�j�����Ӵ�,x=;�Ϭp����L�{�?!1#�3��]���i���d������*�3%i�L�*H�鉿\��(h��W4 	�sK���x�����i��wjQ��[1(�����
�|��7
^U�좥�l$b&`�2�b?��X&��^�:� �(��` �(>��w��yF��_'$f���̟fHĭ�2W�M������K��Nw�ak�n�K� Ax���죑�ر-��R͝�ǵsÚ�*��C�^�$^�#�k@9���s�ڄ6~����S��vM���[EL��8�a����C���K1�e�Lۻ�"��I��^W^"���0�*>�O¹"+�c�P���XoٟF�5vP���5�1�{�V}S� φF�ɦ�o���[It���c��[2	S�)��f�Dt8��M1��
�*���+^ΩO������[4B=Ι
�3>�����R �$W9j%�Jf"~��ΖZ	�J��^�(�B��_|�?�잶�|2,7���y,��GV��!�\�(��LT� �2=�Y����L0��/Ǳ���Ď�eq$07��ADH�!nZ�sF�������������<�mEy�>�]k'��d���1gp�`v껺�6\��>���
k*�HO76s�2�r)����������X�R��v��ֱ!,�'�:&��9�����!Fѩi�푓^H&$9�*4ՀC�/=�\�N�T��*����c@��>N�JzJ�3W�m���ƽ]��Z�T.�g�9<G1`������@N�6�R�fT��LfYJ���i�-�6�hf��^��ZS�*S	�!a4"���y�����U���^��Q�����a���k�gA<�������&�s��q����A��W�Au�x�-��l�����9��B�A��y�� �f�k��VV�]8�)Z��k��n���2C�W���āF�I�EZV���sԽ�T��A�:�'��u�
K�U�O�sP	���h� Y�Qd�ه������3L`�j*4����ב\��b�S��+d�̯V�&)�w�`���72��@�]�=�ç�R飮~���ڙ^�����ޘ��X<E�	���]?��A^.8�$�,�Ђ��[�8J�x���̥bg������Q� �N������J�1X��~��)趁��-y�|7V�� �W�=�7�%�^�BӲ�r%��(�=Ky��$��<|����Y�}�bN:u`����u�J16j�	S]Ш�6<5m�J�&+!��'�3����w8"ל�K4��2�����s�]��
uw��R�+>6��]��TXm;V�D�v�_��'z�/���ZEQ�f���9s���,�i��4�v��6q�M_�]}���<Ҥ�V���0:�Pd�H\#*��27�4iV'���۰�Je4��sQA#�ϰĝ�����lH���PЀs���?$�E���������[�����L2K񶺮�j���Fb�J�]�N�!{�l��BA�Yq�统ez䘃=��������X����ܜ�ɼуCޜ��ir&�s��-�#o͠�$4�������P֔��G=J��oUM_	�EmX�n�l "R�a����YɌ�X��ﯢ�)�=�����9E�����a�ĚF���\_����t����[7���H?��|�S����.��u}ikz�y�e)r��� �S�'���}u]�g@U�	�׬�)%ӝ�PǾ�ˠ�e-Oe@Y!H� Y��7j�p�;_��\�ï�v��NH���];i%�sp�v y^_��wg��j\�W�󁱃��=Î����k!q��J�t!쾙uWМXN��0!�a�2�zMc�c�e�.��
W(,����>|P�˚�2�M,� V	��i9�+4�$?y�obO%��1úy��'��B�2ꪓ�7B]����G��Y(�L��GT�s� ��� qt|A�65@$W����0G��d�3��F�31�+,_���lG2g84�r!)�qYVT
i3b��}l}�B�� �����`7W��GX�����#ʳ(v�O��@9�~��G8ݥ��"r���#�O�ޖ��A��������,4�Q�D^E#!�B��L�-L����x�̂l�ɉ.Ӣ,C�Ġ[�HR%HVO�TG��mj�S�� �)�1��s�Ǫ9�8:Dwt����');��) X(�I�ʹH�5�*��I>Qӱ�4K`��)��BR�K��gV�F1�9��^�~�TE{B�z��cx��\ߺE��$�����sǋ�2O�B�O�'�uY��
�guA���8��I�$?k(�9R�����[��WW�Jv+�%����-��Ƈ�#�������L}2���5����:n(�1���6ح�����u����o�d��Zx���V���u%"c	�]��_z1�w��!�'E*(0["ڋsU��.f/5g�Bj�r���k�����K�>�7̟��{�0�
����c2���34�@6*]���]��Y�����de>��%��������6Zb��\L!�B�6E],S��P�k1]JJ#IZ��%�������UƢo���Y�$h��Z���ϰ�B@������.���풮���֓�>��niR�-�Mρ�%���W�kg�_�W��"�Ȫ�Af�)R�8D�6���l��7Ϧ1j/ɖ��-ꦈ�����wƃ�+Ƅ�rkn���g���z�*��Fw�8��dcE�]sg�&1��y�
,��^��	�^z:�r���߯M�dwu@��@ѿ��6��v�AL�̺�C`��@lɱkA����.��gDנێ�+�m�"I���s�k�*g6�0ԕ��g?U�y�-���Y_z���gP�x(MHDA+����L�:���֓(�~�<�������=���nkԲ��W]����Ƒ�ES�-�ǹ�� ��6��v���o�_ܗ@v��t��E��K"0� �}b�a� d��W�Af��a�qn�V֭�.u }Μ��N��D���(�?^�9dp���H��z��w)fy	?����B���]'�U:�����V��LЪq�kګ�q��ib���)7�>�]K�E�V�GT���܏���b��v9 �Ϥ�x�z��g#�ana�=��#�F�����A��ýp�͐y��-E�ɠ�x�L��������Q':=,��`�H(�g4����G6���U�_�`-Nܒ�%K%��Iƒ�}}�o��qW�^2�S�l��R_D�n����kzo�-�E=��7MC�1�2�}C8�_4z5ֺ��.[~�;*8��/�H��2����F�>�h�;aAt��jbI�y�鿻��mj�)�۵�Y�^T�%^����?�=I����_�!Mх��.�#��*ͳ;+�P<\*t�=M��e�?�k�-����`�M��<���~s�����(	F��Vr�8��]�
N �C#�]J^�N�#�3��m'|�=�����v
X�,^�&���I퉵Q���e��)��o&ɫ؛���ޠ��H�����I���54��/^����ؽ1QOb��z��-���l+�wO�z��вx������c�V�<�����i��:��P����Op���3ɱ������ըx��:$'�%nGe�}�EZ���e�*������q�2�|��azA�_4v�+�9���.0Ĭ_��4>~���g�̃�F���)Ĵk,��Qg���:��V4)�����EUX�ƒ�
���9�>�t:�>�P���m%�{���N��,1��1M�3�{�r�<�x	c+����4z�ut�WJYܕKe�EU�=���h�殞u�F�qb��YM�>fݦB�_��T�=����G�z`F��93��Y��`�� 3�$�)T��5�_�9ܝ$�s���!a4Ո��`ȅ
 ��HIM|��\ l�����E�~r���i�aS�b�g.PY��d�%;G����D�����B$�G��I��F�W�[ *� �a`]�f́V0r�|���^q��w��e��<�חUo����X����s-�'����Iة��?�lB��+Q�ւ'����]��7��\��N�O�����l�뼩B�^��=���ɴ:3���y�ڻf��� ��[;o8�}� /���R�k���tdS�����yjt�iOv�9��7�CQS�f׳!0�&�&��+p>�)A��|R"����-S�U@�|�R�i8"�fe>V��D�֐�[;e�����J��N(ā��/���{M��h.���G��	$�[ٖ������딊��O��D���c���C"F�����o�~���,�S��I�y��15IMM�����4��ٿj�aT i��P/t�}���ر#`r(T���!,���
���9Q��zc��*��6<�Q�T�=s]��� ��q�<��(�$�K�w��ȕ���[���|�e���͐��B�2�GN�CǍK���5��X�����m>ܜ���}�I!s�"D%7V8�p���o����7O�\�e��f�r�,��l�����R�&�-.�"�y3`���f��<�s��4md�K��	��z+(j�+f����k�R�X���'C6��Ru���s�n��r2||wg�f0N���_[�6�`�hV����Oa�Ù�H�7H꾞��e�=aF�O��*��;i�Qh������QvA �_�L��M҉|���T*f�Oٽp׸r�;���zi�|���1���X/onw!;4�li�1	���
���oR<�ȑ�!D�i����T����Y0�NQ�)�>|왮�I�M~tN���m+ �%��&C�x�R�����4[��&7�)��������]9�W�A��)��M��3�J�ɹ�4b/GsbՄ�7��kF��H�̸���x	����Z-�{o�ȈFe���q�����0a��T�`�@������`�WU��=��{��p�Q,���N����"����C>����F�c����7�E˻��j�����uP�d�!;)�a�HV����"Oݬ7=�V��7bnm-�47�Pҏ�V�nf����E�U��D��w�Kqk�)���S��<��m�0��A�׆x<���Ѕ�e�P�ZȨ��t���'Hۢ�B ^���=�<D:��{� :=MfZTҋ*~af�_O��k���̃�p����L=�6}[�]���-q�X9;�5��(���6�x89��l�Mɴ�\<�%���1H�l���~����w	���/�n6�d�a�k`��D��ۓ4��	��9bN�0�m�=�{a�3���vpEa�N`���J3��s�@ۥ44{4P.z-����褾$-��-rjFp5�ʈ�J#�TF�7�o�:H��V��]�(����P� �/��xҐ�K4�d2y��ث��P9+�6�,�m���|�b$����2r�0���`�UXg*���U1�S�μ-- QI\sߴ�ь��7��qr7��
|�*G�V�t!����tah���39^������^��&�+�CS�w��Mcz�`��8�c�ۇ�4^��8����m �h���>��Ɯ�I��̒���ۋ$�DU�����:RҚ��g�B���0&g�r�h�D�lQK'�-{T��G���b�&
���п[�8Cs�&�e_7�����ab�ݬ�� J� �W�Gtހ��uo��|Σb3z5U�0KW)�<��֛DN����9�q�@w�h[�?]��һ2���
���8=֮`�I�S��:ԭ�Za�U��|�*�j�01�B��?�*�#�1)�kj´F��wRi6��v# ��b�<��n�ك�o�T��B����}�EL�:\��A����%n�d1�*���ηh ���b������1_� {ZY~�H~�W��?�;1'�Ξ�,9�ʜ.@Z�0�lJ8}�<lࢎT�,�5��dg�]�ϻFGb/�!��]܊��:��B��j-U������<�[V��o7#�X+e~%Q�̫hW����r�
�-K��O9c���M��*g^hT5ZkΦ-g��*�Px�~q_��z	�	��Nv�Y=��y�Lb	-H��;�Oz��;h�U��D�x����f{&���_%���KJ������`��L�R�)�6��jN؜�!��U�=�x	����j�QcZ6��f
���p��o�ҖA�����5�?a�n���'��yO[j�Ŀ���$$����e�#ė	�
}b4�
K��]���/P2P}��]ʕ:7�`*W]+��D?�'X�{D�ۉg�S 1���R*aY��q����Tp�W��H����?����Ekd?+ǼB�����S��ey�S_)���߻��n�ƙV.o��`ҟ�۬R+Y�c��PN�."��}y<ĭ2��hs�E��� �����&�����Dj	K��z�z=u�V�?�*V#�C!�N$%�Y�*wH��@��=��GB<�_߇p��k\���o�L�1E���-�L���{�o��4��U�p��9���{ʦ����i$!STմ*�IM<��K�E�
�����15�r!|h���kXa:�@Bxd���w�DY�O��=^$J����L'ew�#dd�E��G�km5~��1��S���j�}����4I
��1�:�<� d�e�<e�	#L#w,���~5�R�X���� �9$̌%{���7ث�p}�Z�����g ��;sM��J��J5F�ݧ�E��k�y_i�pf��F������,�q</�)(qV�z�gO��~�c�QBf��)*%οL�^<��%�MM��1�����F��W9+}pJ��n�uƊ��[!�{�Ļ�t�?S��+�+���m3�a�<#��濁��M�~�Q����cBK��}��F1�&'����au�A�F\�!��+�xGX��P�E�� ���ˢ�ύ��1d����{[��~�d��(��y�t*O� �5�l>��X1�0��
�y[��0?����_4�����Ơ���-,�O�c�m6
��xR�Ŝ��/]gIU�l���X���o��,(���/�jK�t��@aV<t���]��]9#1�����6}<�.J�����E�f��>ө.PS,KӮ���S0#A�J.��H3�}K܌���l B���m�����kȿ�`���('���GƠ՘�+������:V�;��N]�D]Ҥ*]^��E�)�qLͪA,<��e�$x�����s�f�	�i��7-��M����I�<;�-,Ɛ��xxZ����=��j��9rW�3��|�'��Y��*{$�t"##:���e��H���~���1c �ól�jЈk���|��q�٫��d}�{��N�) ��ppV#kz�1��槯�}��4��5�U�!����]H4Í�����;��'Um�V5�)k��Hr�.25�ٻG����[B�ДS���[w��9�I�d��0�X�J/�؋{��+�!u1};��Z��b�'o��"pܹ�`G�Ğ�2�ؤB�����J�q���T�&^(�A������\�/����o��
�_����9ܖwd���n�\��`�5�ˬ2���x��,��.��z?e���=��氙� �4��p��¦�zx#�F)�`�gO�W���Z�+Cr
�lK�!�Kh8����%�p��F���W�R��?��C���W��P^��Ct�Ǒ�عTy^�xl�ӎP�^�$̈�?Iם�f0�,5��{�߻��Ǥ��aO]_�nP5'��w\�er��<��TP��.�cܾ�:��Ψq��D8�q��ǝ+�qasExE|�3�o_	�x��i' �1'���"��9���_��i��jΩ!���Y��*(�ٞ~>WҜB�r�C&F�	{tX;������}����5`�<w�^t48���+_�-�sgd~�=�2_Y��k�f6�By�c���7�v���=?C�}���s�qNMݮ�&\B)��	=�A���-_����O�ʦ��@-OB�<�i  -�g�8�ڜB,�dL�����0m.5��VPv����t��V��A�
��� u�������[�b9�\"9�(�x�l��>�A�A[ₐ3K�p���������q@Yd�'�JD�g�o��l�&̡��O�C��ԓek����ac䉁��*M`��^����m��K	���:��%K^`3�����j�摔�p2��1f"F��7&����zi�U�����y�I6��8��V���9�*�%;�FcT�Iy�cW��q��[Ht����d��O~N����f^�9p�����u�>��L���+Ѡ�=��V�VVo��;a;��kq�� �>�>����N�TRz�d�<�2��:�o��5 ǌ�5��S�O�qA�� St1��1®��u^��fJ�	0�jDe㘎r`t�W�Z@�ѽ6�zX��EQ�_���Jq�#V5;֬G�.Q����W~��:��I���]�O�F9Er�z^��m��C��i8���_r�2͐غ�T��9�[6	a\�F���r�2|$�p������Ʒ����G? ��K�Ic�p0{@/���~��81H�wv�~�ȳbz�U��cь�ʺ����4�:��!��SүA"�� ���:��_���Cl�:�7��Ѱ�rWYu����2��66��̩hf5��E)�eL� �&"Gd3�oy�țI}�Z��g�s���^M����d�Rh�fmQ#G�*�����S�t۟b�2�.:�1�d��1C)\n�o_'�4�l�G1q�|6qX��ܵ6�̪-�@=Q/Tߕn5�/�(�Z^	�ާ��<��g�:����<�?���V6�jrMO�]�G��%��G ���|����7^�.��SN�����Xh�^�e�OF1�d�p��x�h��1o�)�eq,��pdew��
X��H�IyD������U�7��K�����[]��*�Ą��'�po@X�i��#����׻�H#oC����Wgd����cWx�V "*a�£y����3�ی'� %�]%��T�9��z����E�:��!��(�l�����e��R`l���������&MN�4E���U��-_�7�O�Q�L���9��
�x��ً���U���"��i�dtĪZM7�����*v����� Լ�VxXFR�A���d,��,��P������A��)�9��b�','�rO�q�@����~�+�`U1���~���Lt͗Y�	�$��`�� �U�R"6�C�H9V;ye,�_84�@Y�L� >��ټ�cv	<�fK�1�^p(�}�[J{��q��c���5\궂�O���-3���W�/��h�Vu�P`Eg:yH���c��%X����(�{��ז���)p��$�`
%�%����8Z/��E�(	X�)���.\�4hI�i����V��y���T��Qퟯ?���'3�=�/����"i�F9�m���b WZ���;	6�a�M�a|2�#ㆲD�H�� ��٬�A��iVz��p�~Me�������LsM�������b�H��R{��v 8����,�OF���ᅊ���i G7�ވ�By�@�Y�r���6o���.'�p�vg*
˼�#[�H$��G�ʬ�[�韰yIk�/�O(���J�I�m���O�~�v9]��E���87<C�rD�>�c���y���9w��E��(���7v�IQ���]�a8s�����ʇ��8�6tq���ߙo'���9#�b	�d��m����/���o:���L�>��Y�͆��S&����cH˄�lY��_ܾW�D�m_J.�Ӓx����+G�	��Rץ�F�`������a6Nx�;��wZ�;J�����\�W��lPG���x+7 ��4
?�5����G4K���H�kLa�u#L�P�-JFb��I�������v��{�XR9h1�=o7�6��ث]�lu,�l추�o���ڦv�P�(F�?x^8�}����Ԏɘ\��%of#��|\����u6�U�z���w�� �)ɀ<�����J1v�R���6}�%ȷ�r��!���Q����jO���Z_M��|���Z0M�B��^�!��w��g� }�D�/�_�5�W���r�7wM5d$$)���dԝnz5jD�s����/1��݃��G���|��W��Y+Jw����<AV�j��]X�DC��Ra={���y$V}SQ�͈Ę������j�ˣ���\��*�{��t�W�e���O�aC�����Qy�fV�~��H����E��VC�	ٻ���
����g;�uѫ ^gy��ੜ`R\�5��n��G
�%���o,�}[��r��賷|�<�r�6������ ܪ�j��5MH�K��AX4�4�RV&r�#jO��hpo].U���Ϙ���{��fp`z]���� �Ѽ��,��hj��b���X�z$&��}:ll'��L��/���q��nUa:bEoF�;�0ۗ]��-c��C�CC�{\�̜R�,3;WC*7t�?k��唵 ����:��	'j*w't`�m���a�=�F��<���l;�Ǚ��N�cc���/hv���5�'tJoR�T�-W��_d�x�	yH�4�c$`�^B��_��,� �Y"���72ʖ�A,��]dSx���	�@����@�[�i���L����ELp�MA�ϲźU4��do���x��Q�q�8�He{G���r�$�Ȭ�0MsJ��|��Q��6��R4�.�w����T?ۛ�y������W���f�Uz�3@�&�en����/[��b,tEV]m�<��Q�����N�t�ݍ"'���4��MD�f�]N��X�^D��8�����i��q3�n�#_��ǁ�##I?����hP�Nm4?b�	0f�DM�����	�X���7����%�:trw�<�lhn{<�3�'w��~�����.ռ�nK�a�/��E�R��w�Y�7w��fP�v�E*�r�%��b�|��q���F�}�
_��
���T>7[G�o"��hpÖ�v�ԝ�i�^��kva��_�^Y1 2�jţP��G&J�΂�Lh�E*GQ��w����_.ʤo���#o�F>,�9��rE��s����Y�o���+�j��i��Gn�/�,jG;�`�&�z�����r�i��~^Ɏ��ˑ�z/�����N~��@7�2P?���C��q?��Yˊ3<"��(nx��SN�d��˗�\� ,��ע�*�̋G��3CLm3�ܓ��Z��K�ڈd��`�(�$<��.�9d�
�k-%�j@3�����5��%	�:�T�#I'��yZ��:�M����T��4��g�FNP0n�u��Ӟ�|�bH.�n�p�"��?f;	����7�3�d9���)Lc����;��u6�e�����G.ǧ`�`vĆQ�3��$�̚(x�Q:�%Z���g�"��o����E�"�7!��`��B`���K<Ҷ�!�@pE6���p�����݃�q�h]46��ٿO�GW�<�`�xbƜ(�,�v�U��Y/;ct=Q�v�~w�28�~P�x_��AD0�|��ύ���ힽ�c��8~�)��Q���ꑱ�B�ԗq&s��M �?i b�Á�˯9Oۺ7@O���
Ʌo���n[Hk5�>P�ɿ��mA�<���^^��!3�m3/==��⏷Q�𠀭"I*�R�y8 �,��ɧ�pr=y��1�����b+�xh�l��&N^�d/���v��zw��=NQ�����Rkwi)��1��J+��L�p�D�5*8~�Ƥ�ˣ����x?~�����M$���b��03�Os�<�ٔ_4��\Gke���Q��55���oK�'�2&Dp���`;e���g�2�bzitRr�����'�~?�e畓l���<�[�D�X��1}�>�T�6훼�c��>`��x�Tl�p�uռ�۠A+I�x���ɶ*\7�N���8�u�w~O���)��������	m�0����V�΄U��Eтu��ߴz�!�����]��l-�?���+�Χ%9���zZN/���̧H^Z	�B���6�_���C���f2�.�P�����YJx+4XP�7�<�DZ�GW،��E�J5c�IJ��V��I���Sǟ3+*2q����x|��{.9r+�D�TXR�x���XyE�$�+�w��P���jo�6W��E��I(;�#r�9&!�ql��+|pԽ"��c����"4X\����D;��%MI*��q�u2
�g!������< ���Z���X�c�fB��{��-V�,	D��o�y3ć���}y�:�d�&@$��[Gn���|{�Q勩fhj�#Y������6>%xY���\��6��4�?���g����p6t]�I}Ie ӵݎ}2BN9�3K��mm��7P��<b��g�G��+֯ �§�VU��.�oe]��������^3�%��-�u0�۫4�����ӗ��iF��D]8�C����]�+��[��c2(7>s��Xc�ӫ��2� �w�3Z�[崣xz������s5c�i�K�g���:T������ա���U@F���<*�!ȃ;%��	�^�ė��b,�W�U��xOسA�C�}4��_���\�����6��82���d�������e�?����V�qq���h����PXGL����o�*#�ev�4����zO�^ ��_"�����2�O�܋�E7Ej��T��y�e|L9T���"'�sS����.&G���;2��%��	�n-0�	�#:�,u��w���]o@\�2h\�$�7�w^Q�5`�O�9���&�BE#F�}�:�����hI#�[�i�=�>�W�Q��e���a*v=�}X��*��H�,P�~7�[�ʦ� �����4��uE�+�Dd9�)Ԓެ�`2h�
�X!��`��МF̖�����E�{��C��I45[�9�w�Qy���sy���*�~�4�l��%��湷�6l0'��|��&lg��OT�⫢�;��k���)��h1�D�.{3����=��-x_]�,4�
�!�\���	K�� �:u}��B�e�i ���N~���Zd.�~dj
(�$��%o{�ذ�!�Y/m�GƯ����Q�^��ab�[&��sY��h<�I#�r]cQ�3ПqO�����ڛ�(#W�"/0c�k��v��qK�01�Й6��+!���R��݈>9�l��gc�2y�6D<,�?;�;�/FlI���A|r�⃊��g���&��3����(m��ָ���B�e|$_�nY7}UϤ|�E���z��4Y�j��h��-h[�{#�*uH�+a�[ni�D��[�0l�?+���+� �`���A�j��H}�P���?�\�rt8�l��O��p�� ���&��5�֓3\T�u0V'��� ՙG�.��?�w�g
y����wT	&׶A2�Id�Jhϱ�� �7�F��n�]��4~R�<G���QRu�o�e���δ.1y���'�qV�Xa4�$�֮���~z����I�i���B���
�"i7�j4_~�L_�R+�z`?j�L�؈��I��Jz��\�s�X�#I�֔C[�f�����p4Bq�N�m<�!P����G&����Cΐ��6w���xB�?%O ��5v��T�/��X�s�mta>��]�<jB0��QDf����U��Du���S�^�����Q�lu�}s7l�}.@�kJ� �"/\�l�"Z�}!�x�j�U=��4EִܜYjzq��O6p0��+��Y��Z�{zV���И3�&l"������k%�
Kg�4�ks^�ao�V�E�1�ekFi��:��R] V��*y7���:�,!�R#Z Ƽ�[��o�M]�k����Á�-&I�'����/!k���q%4?�'[���x�̪����x�sK��F��SY	|�A�<r��j`�
��U�D��f��:��ZY����L_N\tSll�k�C��_��c��z*	ݖ1��jD8��@�fAb�V�5��2�m�}�������-�''��"��g:�v���J��EG��a!*ƥ�Y꽒.�3�QE�]��~v���ÆG=+K��89�q��7�Kz�5�fl�Ǎo>��-0��v�ݟ��~�^��ɕ
{��G@/�G0��Ԭ2��� �}/.B^������<�+�O�)��JgjE 2i`_tֹ捬"6�G���h\�a�;��Ic��(}UR��ͤ�n�h�h��#�q�C��jL#�Oa�S�<s�։�GXܓ�C̅�+�0�By�hc&�,�����g�������L?M ��ׇ�6�1��#S�Hq��o�Ķ.�:b!L���p�em��QP^���_��{5t3���ժ>�{������%�w�؜u�M;�Eݳ���	����C��n�\��9���Ҽ�XY��H�{��+S�߰.��^S��
�J��3/����M���ޤO9;ھ3oL5TG���sA�6�ΨǨJ�����7B�z H��-�i3c���0��u��~�+�û�]#��=lSU�`��W��`� Ou�Tn@�Ԩ�~R:ۘ����ʲ����{�l��Fǐ��Ul��-c�G�y�.r�z������P�2������MN�Y���?�����`����
�t1p�F�<$B�;NhD
�|i�/j���6f�{�<]�Ĕ2�rz��j�-��!�F@�|]! y�Ձֵ�27a$C���;�!ߝ�8Xh����F�Owʱ.����pӲ�};�L��n�MG���,,����@m�}�~��V��'�v�j�N�շ��������l[7�L�����n����2���o����;j���f�lr���ض���&�,���(<���X:��s::�TNQ L\&�Q���Y�U�ůS+�b=��ET�M(�9�#�6{�o �Rk;$��1��a4�O�rP<`�:)^�/�E��@�3s�(-�c@��.�Z��-�������N�e��3��nR~��߯2)p����j�M�I��D~q)��P��&�6��ꗊE�1�4�����[�t�����1Ok.���s��b�Ю4QLOv ��-d�T�X�ܐ����`�ݟ�x�m�g+��BF���W���UX�;mڮ��?�_J�^�Ѧ���Mr-�	B �!a�1��[߀K�V�]6Y�8+37�MX���T�N۱��UR�����s����5����8X�¦S����E^�+f���Z�!g�`æ"�G�W�:C��ɓdbnK�g*���t�tMk�c�o��j4�?��G�q ��#q��;�=�Z�7��WNY&w�vW���ޫ��Աa*�K��Jٸ�J�s#�h�rX�כ�D,�; Uę :�9hj�G,�����- ?0R�h3c�H������?��ͻ~���vu�Z:����L�L�Yv�"
X�r ���+.^}=�v���j������A!?� ���5�O�ܖ9���V�R�}JNs�;{���}sB�ds�uz�<��Բb3�1H��p����.%(Y਽�2�X��4�����<,�#�m�R1Z`R^����Rk�ߨg� 2H�n{`u9#�?�Nî�e�B҄��=o�7"Ƒ�=瀢���(�[u�꾵J�d���s�CS��6��?�򐍇�u�������M�Z�f���������\	�bl���R���$P��3?%�9MyNƏS^����9���^�)?6QC��9N�
`ۙ�<{��69�6gh�.�����V7"Z|[|�ݟamJsL���,F�Ѐ���v�7BL#���9V�vײY�e�C˖�7�v��_�A��h]�.���*h?������/���WM��)5�*5����0[��$�{^�ҧ��
����p�;�}u�	�K Dl���B;�k�[�?Ί�H<��\��E��Uc�C�k�ˬ�!�.�o��;�����t{��0�@��k|28*�i�;n_.�)DԦ2)�j�u�D�K���UU]�{mxZ�;Mw�S�b���v�k�E$<ȸ$���td)y�#��rpx^��*Ďus�P�������˗��$b"ퟤW]o�n�P�6���<�Ы�����Dצ�-�S`�ݤx�S��XN'���sV�['h��YX���.;���O��ģ�G�3<f���#�L�����^v�d�,-�4W3�^qeR[h�}���m��7kNwQ�����Y�p���>�׈4�|�j�EIk|�M�����,G�]�)��;Jw�#A��p�Mv�+�=l�S��՝����f�~f��2�NC��V����p����f����{��c��P�ea��6�3ŷm�7�t�r��D��㻼T�J"<�7b�傊��r=R�+�����jŌ�A��'{�O*�R'�	q�}�n�Ph:ҽ��Eb�e�%�؆ےP�U�[_���U{v��|�\�Y�k0Xjʱ�fT��G��+�ɚ@�f-�]=�+�L�hi�h0������h|Zfq��%���x��5�h�jЃp� ��ӳ��=�t�:NAi�]b����)c[���9/�-�-<2�E�֦v�D�G��s!���7HK���@���V��������Y'4t��l��Q�ki0Xe�Ť��y�l�����zu?��7ILV���.$���2)�;�|T��BM&˪�ݙ_{��cY,9�/K�_��shAH]��rv��'��E�`a�Xb�3����^h�m\'|)��4�kݺv)f���Q�d%t�7���b���z��fP����`Iw� �1�F�#�,����\P2Z�͌d�*ܵ��館�rv���~��C��r6�+��d�U|R�fV> �g��r�a���>��z�	dKݶ)!�@zL�{zbJ�����oN��S��ܙۈ�DH?�)�����W���	��i(NMB���o�����Y.���MV�Atnc�V���Sbş��*��A!
+��	��˩U���ż	Ggxp���c4e����
�څ��_f�e�-�E�,��0�B���)��z�-�1�jI�ZK�a1�j���;��֑tު�L�z���4���|iյ��ױ>4u��0�zn�
�&�z��l]=�T��vz��=N*gkAs{��36O'٭�t�ZR���jR�h������S���ހ�-X;��5NǱQ �;�-}U0"+�c�����6�Y��l ���' 7��)��d�!��8��v�}�;>� �,ˇ���9��aѲ��RP�N�ij|�*p�8f�j�|h�n��
y�ٖW�-s`�m�OM9`W�����;v%�Mu�>�gz0x��gf������z	�D3�oS�"՘���&-HdI��6	X#gr����,@sUI����e�m�28�øn�D\}B���E��^tަ��k�H���D:� 5�5J��[�"�uʜ��GQ`�Y�q0�L��F'���@����=Ѕ�u����Wc���?��Y�g~)z:"պ���,�Q�y�^��.F#��n��6l��S.AR�E�6�����*q�mF�ֱ����tQDiE)�{�@y��J��3/䨾��T�zP��f`��4�+c&����p�|���3>�ߛ�'0�2͇s��:�ݕ�90���!K	������s�������1idP��Pq��ҩˆE�xh�B��j:q^���h���S���A�z�)���`ux/�"F2�p�}���|`O�B���g���VR
��\�%Ұx�'t�� �����,ԵRJ�����+^��jk1�gbL!��;��_gM�w�%]��9/dxcZ��C�p,�FRr��:j��B3fzё*V����elC�����0��Wp�y��β[\KjL""�y��"R��@�L�)��-E��_�;|�z�/j4��b�����;�8"a7ԅ�������uk!�b�x�O,�~V�G&-�a�M0q�M�X��J�PJI5G�?�e�Wh�xu/�������2���4�g8���A[?�$S¶���J%��ॲs�|��n`�[A��k��O!� sϾ��)P�㡝>>Xs�ذ�<?ۓ��D�<��yZ�ܾ�(to�:�uR��beZ�n1�TP@��跐	�G��'����t�2pUtZ�}����#\�pT˂�HG�d䆰ǣ�
��X�:�0V�����w�ܜ��!dN�&ʊR;'�;�f���y��>���j]mF���`s�Slֲ�`1ȗS=��Yr$�=k�9�rvomVζ �!Yqi�C�a��ȢyoÖw�t)���Z�G�9���˻��.��
�Q�8>N���L�G�Y�t#��ݴ�a8���OT�,<ex3�6�svk^�����2�A|�����?c�d�˫��H��~%,� ���
��qi��;��7ǱI���}�B]�
�i2�=��-���~��uX���٬m�)��#ۮ�n�c��I�S��p��N�o�Fp�[�<��k
O�|>N�����h�Hp����m%ֽ8&\ѫ�DE�
	~׿ G,w�؇gB.&A��w�8�h/�xČ�u�ݸڏ���$Qg��5ۄs�o� �������sY�.����~���m��J�{"J���I[go�B�ٕ����9�V(E�3��E�N�;�))�cG=�`ĸ�K�b�~W{E� @�u��,T��`-�B�5j2+�|7��q�*�A�𕰅~+4ʃR��^DdAV��Ց�P�4�/�+���ޗ�(�n��)���|Ph��"�(��R�u�lc�G9��ޝkl�cAw��1�雌у�#	�Z��AZU��7�+�\��[�L+U�ti���Rn�I�ۅG.*h�D�f���4���.>�q6Á	V�n�R44��"�d���!H�;V�nv�¤J�/�}�����:E�CJ�������¼`hg5�y1*��k�����W&���Q�)U[LƖ	�>�-+�FPp߄ת�F��8�=�'m���%qP����)v3v�+��ւ'9�:�R�1-2�{�R��|_�8ٴ�I:��{2��F�*�]�+��,_J��}kKhtk���)$�ǬY���.c_�g��>u���S.�/�.Dy���`B�26�;�,�4s����d�fǗp��t��a�X!��Y_�3�;���u�����Y�n��v�cM!�#@N��Y��6U=ԝ�������ه$��83oĢ�E͘����&��.��i�!��Bo֝� �������c�Y}���T�D Tg� �;E�AA��S�t������=Wff�W�$a�C}=�ǫ�"=��뷅e>Q�Hud1T(c��*Q'q��H� .��l
HF"0S�Tz�"9L�p�j�Zz��y� ���*��xe����N{d��9�f���QX��fy��;v�xӕC��<���f͏&GuM�k�V������*E$���	S
�b>n�n��|���/��G�\$��h��am[!��:u�Z3�ᶘ��!�,��`%_�`�������9�@y�m��p ��8����`���)81���hɯ�8��^@�P�"^LW4�*�`qE�sa)_n�������zq'~�.�s���h+��E�U��U�W���b���:j�w8P��&��+�h��<(9�l=��)J,�HWpZ�Yrb�+`�#	�a��~���	������vB�͖�>fʲB"��������,⋞���v	��)F��{M(���}����[��N�G��2UF�>m�5�פ�p{�$%�NS1��1�&ƘA���)�|5A�ڽdK���#��R��Y�w�F��vNK�"��3$�b��]��,'��8
<15���/������ҥh�K%v	�w�l�\��-y��������w�N��L7AU-ɰ�i��zs ! �t+&�MW�������
f��'��dq�+�	\W8�!A�O�`�z��fCƆ�+E�<Y&8S���x��څ��e���R���֫Q�QA���5�Q;M�L1���#�ws��:��(�>�	�Zr��34k��Q�h'0>M�u��~��m+���;6���1dbsd�3�a�z���ݠ�Nɣ[�=�Ac�OA��g����Q�����sfC���z�%m"aR[��̈Z�
�2r6:�\ثŚe<ުh#'[,���dT��'��8䈣/K���p��!W�bvl�Gn�_��PS�� �i����e�Z.�Yag�����LU�d�N�&���5Fm��o V��t�ƙC�s������	��u���4��IkB�n���EH��)6��Pty\G��*|�xX�T�?�0[����+6��� �����0:��/-r�@��:~���&�������	{���X�����oD� �֡z�xc�<��+g���߃h3p��I��A�Z�P���)�m��.��V��󈥳j�'�^vW�@�@Q��ɭ>��/�f2"��a�~rF���]G^ �S(qö�`I7AH��P]��;�h�z|�#��)�Уa���#���xϿ�Qv`�i~����<OKC�퓚�;���\��)��O��N��R�Sl�$��|��jZ��P:M��'��E�H����
����rɯT����+S�u�����i7#�,��O�'B� �t�W�]�CN�wNG�J�%�O.��������d��ꑓ��.�)�+s08ܳ��u�*���d���!�oB��q�t<^=��|���p$��`��#�����h�<�2�^�$Z�D����S�qj)$L�\w���j�M��k\�ٞ��!!�� �3NO�6V�M�����)�4��!@�'%��O�1�����xz��݈��q�{5,i��XW�kn�
ߞvmS�e�גGr@�]܎������]�g�`PI鶸c���80����#l�fb#Ӓ�GT벨Q�z2�Sc]�n>Po���Wp��ٵ����!��������zbƯ��@�F����ÁU��ڏ-� �W��>+���1B�w����wV��S����[1Wc9-h;�����\�ݟS�p����L�7l���p|'���zD��L����mWq+�$Y�Ս�!�&�犬�-��]/�a�|NRC���Z�,����J���{��ZX �ԗ��w! �|b�|}VD��x, i�v�\��b�jm:�>�T_��%IW�E_�B������O�Q�DGJ[z�H��#�˫���Zu���p�=�#R��D��A _���b���y䍚!
s��x�.Ly���L�s�*�nmpt���d�����~�*A�xġ�e"�1�SPb\��f�w����A�,�ӆF�y��8z蔜�~Ȱ�@�ja���!:�Пe��V�9n}e�I�"�&���X$K@v�'4��F�w�	�/z#b��4j�<��ٻ�<y�7��o�;��7��<�7G�i�V�Г�Wޚ�����H�Y�z��D��h������j�NBgw�@7y���Ϫ������ͅm�mp�5��o�Y=�!��0�A�]9���[]�#f͓����o_�I�J>�� y]�ED�G�Θy(�n+�/��j��r��@��/�51��:�pv���~����'2�u6�@;E@̭��j:x5���%�g�����9Ԙ/en���/vaU��v�	,�֋��-3qc�^yd�MS�#��WA�	Fڄu�l��f�Bh�����*%U�׋��W$��a�pt�k�kc�;ү���д~."��v8��B����bm��ET�YE��e��r�Gt(�QOV.Yj^"��Iz����U���XT�a�)*������jW�Z�{ƽLk�(x���_Nby�Y^I���>�Q����6s�L���˃a4����Zs A��)��qr�kk6�-��@~�JJ�.��OK�JP����fl�%}���VS��/ExY�;�p���X�3�&�r2S�����	����_��ߺ�7ƱL�qnN*��J��٫��$�r������)��o)��Y#�B	W1*Vn���L�*�J�Ā�Ǣ#q���AI�zh�$��1�e�Q6�3<��җ���]���Q=�f��O�!�9�?�S�V;	~' DW����>��U�KY�̅l�����:�SD�>+a��8~�iZ/Lz��i3.�IP5��u�]X�3>o����������>� 'H,R�÷|�D"+��*�6���s���˘�ӜA�Հ��9b��]�P:5��&��W���	�VXt�!��s� Џ9	 I��s0�X�<�d�=g�)I����X+z��)��F!�	��?��#���P�^��T"P�T�.�����3x�Yx�U�޷O|j
̣�c,c\ M�56�[�'��5Hع�@#I�&#ܩ9i����3�����W�^��Cc�C��ܝ�]ԯLy���治�W����{�k_�Ww��v��o�,�ؼ�!��� *�蕎���7�F���sg�B\꼢�Z[�*	�ɫ�	fة:`[���<m�`�8�W��,��)�LDD)�%t�a�
F��Y�Q�w�q�2-b�����f�ʈ�z6lj$KIw}���;��hiϱ:���pF�u�*R��Ʀ��%h�B�t�Ϭ����LH1��,q��p�׫Fl��eE����v�!�ië9�yJ�����5LB+�s�?*�e����,�GY�p�s=�XL�Jql����lGTL&�N\_d�Z,LU��W<߇|Wk?}àFX�!��J�)���0���Vl�c���'�\7�$�EK�vP���X�0�����C"��C%T%�ݦ��\�'rŕ2W�j�9@^�O�fu�<��(�����"c�לCd2iw��y�!胎�nh���G����ˉ�����"i�c���߀+�|�0ri��YC�Z(�Z��5wM=T?�0
��DW�+:�."%�_"�S\k=�U�b7�6_��A�ȟTK	��^Y����.�:n����uT6-��Ə3m��aha;ׂsʊ;���I�Þ{0~�s���z��ҿ���7�����>�:�{�,J���_�;I�ف��u's�s/�!�A>��=s5)˪�L�q�n~Z4�Gm8ݾ9�M)]gX��Q�2�ϭ��N���A �^Xx*��U����&r��!Suީ��n�H��/6xH<�k��Hp�����y��/&����% �#ؾ�&pm��*�i$�ⶱ�0��꥽0=&K�.�"TO���|��Q-E1�"G�������W���XȘIɑnY2
e�������:G{2~˼��p�5�S�"� :���V&��}�CA`��>�ۮ�
��DVǀ�ѹ������1�*6��#��s<���N+�jE�گ��,���O^!��a�qy^'���
Q�a����O�F��~A�ԍ�2"�� ���]p�s5�pv�����i"�0M��^��Ѵ��u���I�����	v;	�Z+�\4�:��B�A�D�ߟkO�@��(��&{YI�(l�, �B0%8*�!��U��1�>��c'�%+a�٪(�I��n�b; vLWw�~i��06f�	^�6^IB͓�Y�����	J�vd�7K{f�W3z�r�-Kb����}>��k���0� ,�*�@�B�@|�W2iA���|�'�q<�J;a��EX�DN�-�>'���;�_ޞ��|����۴����Ws�����"��4�����R�o��eP��D�׈��E�]�s��vX��=X�YKr}�Z秢1u�h}r}ay�f	���f0|n7mϥa���*���`�-�,~u2����)���B�$:����!��^@�"+��X�S^Z���>W����|�G��������u�;P�".���^�}IK��}}��kō#�3�����5�u��>8o�����+0WFvEm�=����X��Bp��}!�g���oU�� 
g�92��kk!d�2���In����>�UJ~d$��
�?)T�r�u��ǉv��Cb�o�A���3�	�D�h�%���.J��FRѲ���2����OW,y�k�ң4u�>gB?~��]=L��É��Y%B�}y�1��I�l?�b���z��#�h�}���qV��M<P>�E�f�$C���3�"rq�i��y��3#M���ϒ��,�=�}��Ilji�i�m�oyS��NMp�c�ji}����n}%Ji��}����W>��^��^����Ĵ�
�m��Cb��3���ً��6��ۘ|�,D�^��*T���qW��	�'�d�����Q6C~�jw��Y��a���cXAv[2|0��-d.*�[��{����_/����a�a�Rk�X	��d�p3N��<�x*O�w~KET�RdVy��_�(q�ss�������h ����
�g�Nj��g��|'�x�̢�F~_�apR͂������l�ct�m���&]68<'?�ޟ�l�@QN�����ǁIT�)�i�/�uR��@��:�2�>���]��TJ���QA \�~��Ñ�8Ckj*�I:�' ]�	�Crc�L���r�oYo�j}��u�8�'i�%���m`�4`|�����7�9���������:��I��v��>AE�5'��{���=\G9-,B����}�,~�uܥ9+�C��Q�:��L��{�����rZ�<]��IS#u�Z�>
p �a�g���#��b��3�
9��5[|m��BƬc, �&��|&0�Y�o���(�<X���ȝo�N�Ï��@�CLt�D�[����m�Z�~'8�TX����#[�¦UC�<�[ҔaP�~4�3iL�e��Hc������Z1n�R����>�d��;zdZ���r��r�KbI#�"bC$3xh'�-	����0����V��0A{�`jG�9n&S� d�[�;Pq�s�/Lg��xi3�����uD+<�F`��@�ܢ�_ё!49�-���ܑ�?NJ㇙�u��[,�Y��f'�)�>�����|F�"Λ��/?�|?��܃-hzD�Gn�,[-�{;� �`@�ztZ��
A�?g���Y+�rf�o�Pw^�������I���x="�����'�1ܓ%�7��n"��7��r� ��C�IڳN����\�k���M��e�d�"TI~�\��!�ǖ�c�ڣ#�t�֖f����p}f�y�U��7�y��'س��0�̷�����IO\ ���Q�
�.��G��$�4@�p@�2���9�o�d�[�5�pM
*!0��Z�žb9ש�0	���KVc~�/�M�ڇ��C���$������& �0r�P�?wrސ]<1���d��SEs7jd�[SZG$}�e%]u.#�8� u��+v�sH����7��c���
�>���/�Ӽ�6��3*)�x�V���ݔVD�\�:&P"l���|Ht���e<o��
�4O���֥�pf��ϣ�qxZ��s��n�*cZ�f�s�=��ht����w���������"S:����S���x�{	�~A1��v*L�3��9�+�u�H⎓a<^��b鑗>ʆ҄3�)#��?�䊥��UG��7� Z{#Y�7��@X�ۼ�}౹^�ë��	a���������޼'������s_m]%��3�u*﵋Oԫ.��"T�R�t9P@]{�w�������"�W,q�^�`��7���`�ӄ}�s����zsA�j��l{�U���f�t^1)p(��A3��I�,H|�J#e'�
�:�}̾��j^� -��M-m��D��"��$MF���[R���<��b��H')��]F�`�s���ӧ9�P9E����qf�nx�sW�m��KT�o9���}.�D?���i��Y>tl��[(�4lĥ�;�.c�w3Z��b�h?�qJW���W.��D�Ć.��@+�Q2VY+���i`vV�D��2���q?t��Q�K�����J/�t5V_��Q��fohY��N�p\"+�g��L͏�v|�\�J%6���h��3ґ���XzʜJ��c�f���d9 &�I��2�=���M��G������w�	�W��r�.��~kG� ��	�\qN$RG��WY�;I9IQѻ�I��w�:|eəUx��Q<?���39���wAV+��A�i7��6�s��J3�����b��Re�f�6�km>Z��Wg��Mw�ZBj���M,v힝��c��,��X��֭��!K�RY��"�@æ+j��l��r͉�:�0��I��4��Ցa��P�y�$ɐ�Z���dA�u��-�e��0����A�|б]���Н�a�� ��>�������0B��H�oWY�_��639*�G-�	��<X�O�����S�mױ�E��;�Ҟ�`��F����Deuع�x��/nz��E1%��� ��?W4��#{����$p����__1H� ���\������t}������W��w������X�����]�3������,uךze���glw��[*��)�ȇ,�d���D#T���jd�S�������r\ω]ò����ѵb�ѡ�:` ����g��d���Hs�-�����5C�m0T<��D"�+�va�0Y�<��*@�g�	�XWb<�m�l�amsu�[��7j�6�'uc�Mch.z
r���P��RYU�]D�G��7VZOO�^��e��oi�p���3��0MI>L���[��L���=_�ܝ�f��(N|�R!��CT��@59{(�xH���il�`
I���)ݢo@~)o��S��1#�1���?v�3��X�� �r��Ͱ{`�wN�Xdy������DX�v}i�ͮ^i� ��W���n��rJ�! z����Lec����J�#��	
x�z�₯���N1���<O�aw��U�lo2�mS�����)��=g���Zek�٨��J�3�j��޲����H��װ��;��lA�ky�
;�u���lqt��y�M���E��#��@_u��1+�1ПZ�
��~:|�x�I	6���$!k�#���GN�L�!��"8��n����ad����F�&$J@��DdA�8K����I�j�wO@�3e~&��$�b��&1U��O?����~��l��Fä횯��I?ʳ��MYu���rL��h���y�%�e|�ӷA�����勷������T�t§-�����(���^�y|U�{��#W��,<��50QD:�d���D)e�"�����=��"���6�4F����0��zT�9��&�\�L�@}����,x��0���?Q,�/��+�����h�~4@
g�s��PM��d�-�-b!���5����C��ܦ�2HZ��v��`
�m��V����:��}˞�LO��A}O,M�7R�1{Q2�`|�k���͈�a��x��tK�";8�~N��>y�~�i2T{WL(�@�p��&��U���o�(X�?U�� ]�,*a�J����e�Yc�=1�����
E*}�4���R�˘\]�Mr���>�X��i�(��x�9�*�H�N�������ߣ@5T����.\r����������Vu]�?T/��b�@i�_��$,vs���M�!��~N���p!�o6%���т��^��fLD�I�]_ �-��r"O���?�3�ѓM�CI���*�G�f����9V���W���\N΁�Yʗb��vG0���g֔�lnB�k8RO�_�ˢ�(�"�4�tS& 9��)D��r����]�+91zdݼ���JNZ[��5J�J��!�:��R��u���\��*��������P�3&�ϧm�w鎫g��w�7��ކ�P�%�g���䜰���Xj1��t댺]��4��f5)�H#W���b�BCр���Z��-�*M���7��l��'��7�Nb�W�C?��Yj��������YR5;%�޾���I�?�)֌3�z'ul\˳g�,B]�*��g?�N4!�a�"6����<f.o����!��s�x�6Ѱ��p���c��@��j�!a��*�bS�~<EN5;�������
�� B3#C��V/V����|���I��rU�s�6|���E8*r����βJ��+�u�p�*a�.���cZ�����O����O��"[TiCc3��]^}�d�Y�=[_��9%��1!.��A�uC�g'>�YD{��r�{Tؽ�j<�>���Uc�N�����jP��uk���(���� �j�y��f3o�lr�]R�h(%�P�
�ۻ�l�i]��Y�r�B�z����=���n��Y�=# �i��O��ʏ㾿����$����?_Wʢ<���m��)l��23�g�?�7�}e�N_�w�w@�]�V�p#����[ED$+�Q
7�C
!�i���6u��dv�k��q�c*��I��6oY�'{Ҥ�j��t����ҭ0!çzS-7ݍ�m�k��I%���vK��.4l�2
ÿ���Ixa��\R��L��ջ	&�x���:,�Ϣ��e���;]æ��R[�]!�W̰�}��ɒ�x�U�-?����}��M�p����>�$?N�!�.��KpY�����VH�a�=k�]͹Ԏ	��W�]%^;�`L;\�|��Č+�Æ�m/yO��њ8���&�ÑN	�tkk۪D@�����B�ʑ�L�~��j��a�Y�Ŗ#Ke/]�@�`�گ��noJ��+k�R�W9v0��������~���m3��+)�� @=�P�Wk�D����$��;�s��|{.��6�d��q�ET�9{kC..]I��p���M+Xw��E�B��p��M�Mʺ�a�ԌF�(kU��S��Nր5T�Z�r������W0�xV�M��պ�s��ELW��xjhp/
(�R6}ɜ�I�T�c������5k0^�%x�F��EeIC��h�B�0ɋBg���X�l��.�(���Cέ�'�(���q�y��<��z+6oոQ��61�N*�Q5ߦV�|'��������p*Cz[�ѩ�m�?���Z������厷y�	a�TT�������J!�Jx'M}�� ����Y5���A��"�Q�����  �,�����>X��h�O���[0���Z*��,����R�����j(#�r4m�qZ��A�^Xis��%���V����ʳR��3�H��Z�/�BYN����_��]�S�b13����:��Pz��D�;0UWĒA�t$�n#'��7O�)D�K��n�9:�bk>�`��/D��/�U�+허L-A��e�᫏�ǌ��J�J�����!��	J��T����LX�gO��]	u j��tv%"��� ee�ڗ$Цy,�*g�,')B�9�sχ��4�o'UqGa*�%hΫ�5�d:����}_��-�J�~h�KC���a��ؒ��XX�6�HtI`0ݝc�>�N���l�B���ҫ��-�_|Z69'���Rw�C�q)Dx�����3g�CU�����<��P����~=I>ׁ������Q��_+6w�ѝsgɦ��(�nT�f��Cl|��@�X`LxeJ�b�ay��Yf��s����p��vhG���p(�W;���0�
h4m�,�)�Y���W��,�#��	t�1�P�G�G〿�!�����R�m�$�xZh�q϶J�8kYcE �M	t���H��D�-��F}=��Fx��6�n�W����G����M�(�'"�#@\�	�2 ��Rc�:�^��Ѽ�*���]%��̈����L2�veO�6B���$��3vW�{m|�uw[�-�YX�'r,#�V������P�l�j�T��	D[!�h��^0SNex}Gɫ�\o�e4ٿ
����P lɷg����P�i}�2*%-��%_�Ėq�g�J�_��L�E��tAӀ����
�����q�@�VzB�����\��Rxy�f������voE;k��2����4�MRM��9����n$:��6��{!�����Q�X�q#3WT��F�~�{r&8�8�R��O�_��=�Q<(<L��Jc6m47	E��ҡ���9!:֠߯���a����(�y̲�?b\��ҭ8Aٟ)G_?e���.��ђ�<��t��.iGY�H�y�dSm7���{V39�T��t��R{YkL��@�%�a,��up���[;�i�����I�m�8;v:vʒ�Rk��
����I�Q��*,v�����\��H���>Ze�ѹW��D��P���m\���u���4e�G��a�'sP�t�@6�!>q&������p_%�J� d�q����"2�e�JL ����$[yD� ,�������C�O���b�p� �kk�9P@��Rɒ���"�a&�q��I4#���[����	,�.t�mH����O;�`fs��ӂ!�˵  ��F����4�a��څ��mb$��-xU4J|�J���=���Z��^���R�*F25�gKj־���Վ[&����e��ƢU�!_bA6�p}&��۷(��H1���rޗ0�ش$�Q<6���M~��Y+[�2:�v�s�H�'lOMq"�S��[d|��\�����By�	V�C�j�����,�gD��h3�zH��q����<��3#I.�$��.[��j�Z��G	�����p�H��Ё4cb�¹v#�����jxR��vR��y�6��
vǣ��q������7�@��n��-M=B�WT��|��u7�oa�g7xH����؅�|�Zy'�{F���wa�?������]���݉��;s5�̹�P����t��'+[^u��3��3@|�YB$�j�����.-��r���Lq%���S �������*�v�X�̾
��Kr֥V�(���
ǯIR��*�)��D�I�<���ܹ ��B��j1��TD�x��v�8#Xk��r�ͻ0J�q�v�UG�	2'
c|��.]�#!���Ŀ�֖�Ĳ��K�MKhbr�}��p�@�:���{es��5��+���XY=M��ϖ.Y�Ti��p��4;o����!�A�$�~^��r(+���X�r#5�(fsC%Lo��>����_��B����~��jQ�����s��͉bB~+�ک�tIc� �W��Ad��?���1�8�:A��|)�"y�z��U�]GF ��a	�E3�hL	��֟I��H}�FS4=�d�8*���i�(�`d�zކS��ozxS��7�[�=+N�4���>M�%U��`�PW�
��!xsF8tI˝D��3���$�,Y	#=W��E"�9�ć�dK��M���bT�i]Q�
�V�}X���g�'j3(�;�t�������<�J�h�����HP�T�7�����c�3ʋ/�Md���3/E�
��8Ӿ���?b�sJG��T��4a�q�N"�E=7����^��&ų�Dos��3Lcq�ٓ�m�Vr��=�T8ɟ}��1Nks��2Hǁ��_h����#ZX� �d�Z׋�7�F�:˝����(���ϒu������T|=F2�Z`XD�)���
M��>wp�6j�s}3 �ku3w�Z,=Q��ˇQc�s�\�#���6N��2h�B�]��LzQs<�P���FH�e�g������"��pvK86J'1ί)�v�-����ɫX{C=|ĉM�0�(��Cg���j+����$]C%iϽ���p�]��%�@+���=y5e!-���߉����xv�Z%r�Yғ��NZß�<̭'u�")cqo:,�@��J�Zs���g>G|lF<q���sA��tp���DlkE�h���ڌ�T�L��n1�@���ƀ�ڤ���H�i�o
"�k�^LG�X�6�X��z\�@j�*��R�Ęr�3D����g����T��Og{0f#��p�?uӘ�r����'�E���cވ-h�Y��Z�4<��`Xu�e�Hcp����m����"��~ό�#r9.��̱�`[7�A<�p�p��*񾃰�]��GT�/�a���U�s�o�*V+��.[O��[M�����֬� �L>��yZ8����3"nT�|f祈��\gzU�5接5w���'hPћv��2�Яb��3��#�:Oճ���]ҕ��|�{��v�}�ķ�Ų���kF�#�����<�$�r���ӏ�4a|�~�-l��fXi1�O�H=.�
A:#��ƻ0A|v5�)�����JtJ�S %�z��o|�kz�\^
��Z���u
��?��H]��ei��Y7\&�_Xp_���r�����ptr�>�}i�tYg�R@k���u�"i<|vB�K�b]Ǆ��k���V�1�Z�F&��'F��y[�� �=���3�^�h���Ԛ�9��c<a�����]�ʾ��q=ڿ��z�2���j(�����-�x.���!V�\�RR�G�M��|���-b�����B������J�ԟ\!�j���m����|_4b`�y2R�Fe��$!���>ۜ&&bY�֤����h9L�g��(,9r��q�.7�?�:7��8K�gYk���-A��-�d��8�0�m��Ȼ�m���g�L�އtA+�<L$a@�7A��v��|��U���c����)�!�Up��@i��A�q!K���i,*a��!%G�L<яr��!N#�ȗb����Ƨ,3��i�(���� T�8 `s��ؔ|Ã�/�(oDIaK�"�Cu^�0��<$���q�>Ÿ�/��L�_/�g�ڿ�y� ԀO����,�&��^x�'�L������M9f|\S�����"O�ѩ;� x��*���1aƒ��_��6��X���L�}h�����ĸ�Ce�D�u₉�n��e��&᠉�̜���)����Ӱ;|8�T3�*{̿Kz+?�U3����d^w#K@��ï!��~���ѱ۳�(�B�u�ψ̋�k���������.�E_�5���5X���sr����2�HJ)�q��+4��D��kDH|�`/��v�*ښ,O��E �_TA��fUcA�%���%'��	h���h;l�:����Ԓ���G��ёD�����
l(�:"��2lrf�q��-��E��{�F�k�>IQ�E�=���<���Y�*}x�Q���!����l1'�V��Q���3$��SQ�=괓o�
��yG��`tD�Q���a�1K�o1)-Hˇt�8�H�n�R�Ȅ x_�V�/z�#�_�ֽ����&������5[���T �Wp ���Mw	�i�A2��=���J�a�ڵDL�ξ��|���C����c�nᅨ�69�������qrV3�Mr࿏��S�^
�.���8�cGDg�J,R��d�����U�zW4�]����ʆ9e����GXT�n�8t v��[M��c� M��ڤH|2f�k���R31Q��|l����+h7���k4?:����?��{#k��5c�N�G�|X��5Ս���$���oR��ꬱC�
(����,�(��].Q���@�W��C�Pi����;I�r�[�zN��Q�;Jbh����ʻ�d���������5X�j�ؐyq�f��0�XW���m4�E���Fۢd$�!ަ��;����z�]�
<v����~���SԐ
[�_I����b��|�d�j�W�<�;f�CM��EGq�YT�w��)y�,�AO�xڐ1�����'�9��\I*� +j��JMi�a��D����D�j��m��ѷ_ma$z�ӗ9�P����4��G�o١��PHy�K�/8F��^H40��K�N�E�,���˔	eF&�`�'�\� �{ė�>Ͱv���J���P~SC6���?v��+�֢��U�*d�.o���Xˤ[���.�n+���|U]Ԫ��X2n,w�9s+<����,5��n^o}��TN <�"kM4B�U?�}�����$DDжa�BZj����Y��rj�gZb!��+$�Vx��������m����1d�Oq#�2Q�/��^�jq�^�Ȥ0o.�V�8a���?*�y]�b���u�ѹr��U��S;>��@�KrQ�c�\Z����B��Dx R6��nñv ¿M�o�i1��\�|A�A��Y�4 �{�S��E��:�J[����r��;�~8��ߙw�8��?ّ$�v׉m�;l���V죸�Xܮ+���v�Fl�g����>G@�+���;+q4�^
��l�a��\��.���+�[P%���Vd�Tv��!*>Iӳc8�I�g� �s���@Q!l2��������Nj��GT0^�����[��4?kS��3p�v��:�i�2G�\��_��I�v[����p�0,���l,�c�p#��_ �A���x�^]]Ɇ�QT���N�=?�㒼 �8�P��ۢ,�"\�Q���b��TFH��� c1&1PF���ρٛ�,F�u���@5�CS%�q�thTʺ�����u`e�f�2��n���iɒ K_�	������)��E{�x��^V;���5`,�?NeV����	�r�3�-%0�G1�)�u���l�������J^�Q,i6��F�@�caI�x_d��N;;*����CM�y�9��o��OE/@/�<˙����G���}�%���Cw�F�����*�܁���+P�Xf���>r�����_Wȫ-.�	�	��&gU�:��Ub��u�h~��s%o��\L�Y�9�rљR�
)P�s�w��E���GM�A<��z�|�L�!@��"$��K	c�8�g�U�|�Hc�!"��(�~9��_�炮��m���$�e�Лw�lw���_�!���2w���3���ݍ}f#��DL�0~dפ^��GT���\%��~�k7"ƚXse�2�q�!~T,_Q(�x��bkWm�q�m]s+l斮�z�!�y2��ohZ�F$X���ቆb��pu����΄�L�gy�wû���. t�L�]8L��-Ƣ}Z(;M~������TǱ�1$��|kBP���`�����+M�L�  +��1_;��N�g]�T����:��������!���{S� �i�n7'���� @y1��lOo���m�o+i�pL?���	���\ʦ����X�|P�C]-{��kIH$X@|JO`b�6uPOz��4"���P�a���4C�
i�~��V�u���䱂��}�ץ{�4����n6���$<��}1�FB�*�-$ k��Ax<�k�;����=C��z���02��$��]�q	����N�k6�y�FcͿ���	u�F��D$,3W�B�\2����R�#l8�ʣ�����\����au`��9���ǃ<��lJ`�L��K C5���.��센u�v�`�Zyc9+�7Aը>#���]�>�K�r����"z�$�o�vߝ�T�SZ�ycM����PܱJv���<_�%]N,�'o	�Un�u�`����/�ޝc�tg<���X�P�%
������ޯv�4�+�bDF"CE�F΍��/{#f�|GE�;9��QS�����~�����.n|�,�I�h$�QJ65D>+����VY���Z�v���'��#�Q<{#���������K����	�N<��T}�08�p>G.�u��"���=o�:�:&-�	����.mϐ�L�-?�6H�P��������G��@�&��o���hEg$��֗�X�",�6
~U�̵�}|���O�t�ka�h����w���*f8bzÍ��M���aS7���B		��J��I�u�~� �!%���o4��VG x����K�\���x��zs�w������D�q�i�������^��օU��W��N\Px�xZP>qku6�(uE�e3E���u�������Q�|j�M��#~=��9�X߉B�?T�&ʋ�B@����7��+�5�Q�3��7�d4��(��Z79y�yR	��>x�Gi&K�g��A/*��mQ�u��5o�M�F�p��(D��e���4���>N�Z
ɋX�5�)���H�xT[�a�zͨ�+�Z��9��Ղ�*m�a�j^8�/5;��<�k�˰��DOsi�>�_@r�S��(���*4��5�D$M�=ޤ���v���_�؊k�i�{u�@�4n��T�g���-M��u�":,"��,&�5��(���8l�}n�^�1��Nd+�����%e��{�]8TKH|�c�Hʽܜ���1�{�8j�iZ3�U�ɽK��Ɂ��E���/��WԹ��,)�P�G�e�����\m�b
�ъ �Q�+�ƪ(9�P]�iC�<���a��� b%��& ���r���I�7��%+)i�)�{E���|����s(�`f��dZ'��6�8�B��<K�%�Q�$/��_���/���շS�e��`��ZHa�콒�%s��_d�
b�ch�U�1��hF��
��Fwٷ �e�\KL������mڍo-7��Xh37��?:��F�G؍حV�j�	[qcM=I�v��1O�^��) 'n����Z������y�O���R�s�n���b��js�g������3V[T��V����*���̆�?8E���1ܖ�E}��1f��?��n�SHB��#�Z��<��ŰP/)S�0/�-Qo_R:H���nMm�-xc�wovA)ۜ�B�ڲ&��0o��]Yg��]�p�E�V�mA��1m��E�q�v�h~�q�ɉ�쮎�R���o&����鸑C�j�����涧���|ɛFZ5;tЅ?�zf�fm�M�	"7�w$/�D; �/k�y�O텢�Oh���੖f��-�����{R*{4jבs�T���m��&�C���_Ko�(f��rz���1c����1V�3䥽;�85@�����SwJbzvcM��2߂��Du�&���wB�������NG�� q~A3%>��.�x��K3����;%�H���6Z+�u�z�ۨ��hrTI�dmď����95i��4e��%#,Մݫ�z�7���$񱷺,k^Qzy	͋bq�T�
jɘ�U]��HK@�w��,q�i-��ZU�!cs@��Q_1���-5�;�A��S�VM*���-A��|h�.4�^�$��n[��� Ǉ����L��שy���&������h�	i2�뀎�W$�g$��F��s�+q�e)�P�� l��j�q�l���{��1��ܠ٧�BP��?)�Bɞ�常Ԑ32�2r�y�i�ԢţfbfzM�JX9?�4��>"�P���u6��j��m;��J�*z����������C�
H���^�3}#�b����Uk/t
���/��`Ԉ������IJp�2^|�����O˒��vC��� �����V�V�VD�^?�����vM �^�BNH׷��5k��=9/² ��,�m�%n��u��AN�V#�������p����(��Zd`����R�<���|3�zc�3�P���~�'/]�������մv+�r)e����ÇS�W��\7��M�57�Mv?T�?�JJ��˞�n�8�r@��x�����A���͊(��C�ѳV��q>8C��"�	/ض�Q)��WWs����L�H�)��ߛ���hӛ���{�x�����q�J�)�޻�Ijc����~�g�A;���/���ZTv�Q��.2f�d�S����~�=.���QЧ�#B~�Z�/�ZE���Kຢ���X���G��Bl	�$�`,��ӝ�1��\��DƄ��v�(r!��*6K�~��3��0rpR�v�Ɠ�u���7���=Wrk�[�![�Q�,�*n>
����+���+e��8��>D�fHʣ#M��❡pU t�˄/sCX�<�d� ipklդ�y��
��+�b��e�l��C�f��z`x��ҙ�z��	%q��JkTh_�uW��� 0-_]��k�ͥ�@Y=u�OꘝehQZ{���rs��\/H�C��~��ik�4���1~YSw��P���i�����"B���ɜ�Y�?�� �a�xL@�aRp��T��)�����u_OH R��BXT`C�7�3*x2epz���N���;�=���������	�w�Z��T��1p�ϩIi	��{g�34�3�{�M�m2�n��߹h	�z^4ЛD$6	}�|�Ҙ�R�RIy
(p���)�}��$j�8/F-oDq��삘eۘA��٤B��
PG�2WpE44���/h�]~im�˥L�����š�6|�e���zZ�З�'s��)�kW� }��+�X��7{`o���t��yq��m$PUj�'$�+Yi�ӵ�����,��84��"��aXbK��W�b��h8N�?�:w߇�%x����j���yfص�$�0����_�� �(��2����.^��_�hPA[~b�L��Q,m�v�p�c|6ީY��{�e³n�u��wI��tv��ϔ��%�r��ryJ������
cr�Ϭ*Y>a��[M��·ٴx�576ꘌ?w@H�s�m�W6�����.\�Dy�t�fI��DP��(:<}���34�sf�
��J��z'��d��L�s��p�%�BqV�o�t����O����-�Mx�����$���Xs�� �d��S'P{y�}� d��&����wU�����O<�<m�[L�%��Y ����/����]�R�w#}R�}j�<��.�̞��}6�AA���=u�|~C�\x�G�'�3�8u�q���'I��f6��Y8�ZD'h���g�MDh-�Y��m��*	7��7��m�Q�j���e�Qј�u�U�2o���b7ЂJ���}Jrm��R�,I�U!�'��Uu:�S���5���lB0zf��7�a��;�E�B��ԉ�𐊊#�9;PhH�Hr���� �lỴ�[u�	��h�Y���&�f�����K6�/<#h�>U� ���k�m��Q~�
m��!{g�xӽ�bF�[���R6��IP��9��� �Ҩh���y��P�z���A���0��>*�l��Lo� ���"� Q�R�j��z
/��
�;f��y�#Q�C �AX4�����<or��='��eU7^�����T�o�C�r����}/NW-��%ǀժ�����w��ޭ�n}�G+x���{�_�t_���� ��~����®2����x�	��r�^�$0#�׾$��.2GXO�)�w�L�~y?��-o���W���+��_w�~���F]��sa	ED[�B��f�&�i/㲑���*��GX�(�y;V��;u2�9�Żh1��lOS�}�}iԨ���z�+gx�f`����7��R+��<o�Z�n]{݊�����s���\�P�c%Z��$-�%��i��*G�7ٿ��ŏ}�Т�N����8Z�T��~��`<٥��0K��Cx�c��w��4�9Nɪ��k�W���q@a ʩ�]z��~/��(j�U^2n=�w�{\��1&-�0�wGo�C�k��9<��9����,�D�mK��'�n(a�	���{C�x�(�}�m {�C���-�l����؈��3P�M�co;�f�2eQxʗxe�eV��@�68E������!�ȊW_/7K,����t��1�0�~f.d�m���ꦹK���=x6UNه�,�o�A�-�q�_���K�ެBO�!Nk�)'���ǽ����V�)B
 �#U/���g�]�����타@�|(e&G��&v��6<�qǷ�>;Q�?��tN�?*W��%���UzBI?��ݬ�yUwF!L���;�!!pi�2�{2�C�֠������L�;��Ҭĳq��J$O_cpd][Ϡ&f��i6�1�@����O(�T�N+�z�Y�&�Z|*̶�o���E�_+��J�K�,:��Q�:�/����>��q2�c�<�^˒o�"k�{cB����	ƛRJ��B^�J ��P�^A6�j�2Z�%�tcg�ɍD���V�\��0�S�����;d@&]���UE��:Q�uZJ��R�d7촨�������G�C5uNMχ��(�b$C?I��i(ju%��U|{�;z5���D�K�W�r�:' �M�)����d��X��qa�hhi�ػ�p��_�ܧW�~�[���A�ܗ��dْ�^)
��0�L'x���y�r��5`��DܱO��ֶ�y�,�u���E�7�O����A?���Q��^z��5hJg��!��嬇��g�*d��'��bO�t�S\�[�:-�ô�ҽ_w�H3�=�k�̞s�BjW�zI�(#�pw�8`�xH�����X��GQ���W3�.�h��A���\Y��N����J�\�DA{-"��f�ȫf,�-F?�=�ヒ�2�rj�M������hH�)WT8��\KX��9�<���aբ�	��>?�o� ��a.~<)3�� [1�s91Oh� $� ��:�8��iF�{��Y��S����9~g@���|F�������.����Cjn^gk߮��+@K��Ü�E�p	�fF�$#�m�q�����Xi-�)3/_r����夆�I#h�W���>��S��{z 
@�1�h��I�����6O
��&��"u��_Jڊ`<�p9^G�4<|�Jxblx���3t���oac�����HqK��?����c6��F�4�Z���=�M�&!�W����4Hkw;(��0�Q�7;�4Y���pC��*X�n_�-]��A×:'e��XD���,�n�?@�J������Y�&y]�S^��D�wX��,�}yjχ��Z���F}� ��L#��e��HH�%��p7;9F�:�3ayO��#�*6���Ԕ �������û�q��9[�6�0���gQ��Q���𗈁��94^7�

���v�2#!��.D�}YϘBor�,��4T��y�$嚆��	���EU�l�t#2a��SJ �Bqf2���{�qg��;g�ɤ���h�� ���3vzz�ҫ�Kc30J�Bl�<����$?�>/dH���+~�toװ� g�j`,|�շ@3��6��	����-���r�^R�d�I3���Ei�]�U��k�g5�sN�h .��f��#�0�n�r��p�lwW��*'[�:�t��@ �O��e'��R=g��{c���
�A����{*�ݦ��!Yn�?���s�Z�g���z�n�}ȹCk9N�>L�z�q-�db�MM�I��&�wb���1J'wim.�*���j ��]�t�JME�q@���yU��l�:���7��c�' ��
ڄ	$"Y����O�rlF��&�e�[�te��6��6{m/]��a�L�٨e��2�sr��!��/��e���z�Q��y^>���|��@*ҟ�t���������M!G9�Z���:g�y������{�|����
o�SΌ�uC�`Q�����S�l=U	s_c&�w "��2��{���~q��ç��9!��w�Qq �
�9�V4}�#��/R^_<�Ξ�0|&������3��@-�.U?I��Xiw�Lj@�8Y�Nr�sܐ�jn�SG%\�-�C��X�h)��@D2��n�hx����zw���$�Cޙr�@�݁Y�Nc�=��!A� ��.��l�M�e5X���ja��h'��+JCI��f:S�ȀL�m7��m����u�FI@T�U�[��]VkB	�N;�$C���Y�?5Lψ��ri�C^3��c4}��VTw@A��� �V�Zj�yw Ǔc�7�^��;�����7�Fq����^�4��oa^܁E�vc�}��7ڼ5d���Ɇ@��+,|#��9�2�_~�R͊х�3�ԑ~����[����`5
j.���1m��"#��j��5�,�'�����g{�~~�
�i��֧��:�MN�'yV��	���4���#A�2�$�ս%t��dO�Tjp�sL��I�
�V��M�u�
�&�����r/i�~s�B�c���J��-�Qě��w�q�c��	1Q�9�,T���7Da�M��Ej���</�Y/.�j�����&�%.e�C�o�k�x��?`�{��柊f�2n�W�~V���-b�Uw�>o�.�e6��5l��� "u��ֿ�B}�\���}�P>���N��$~
wX�>������&P9|�0hAƀMC���*4*J�:��u$�;e��p��q����M��i|��ed���Ҏ���xX�ފ2�0���:�X=*�U�8���Y�GI�c�<���o�F}9����@;]�F��vD�Q
��ї'e�y}���;���1�'�vQ�4��߬4�P��r���t�s݋�	'%����kN>��9����	@1����������I6��2�G\S킈d��^%��-����Ҟ��E��ȡ�V��[$M��9�D ����#���ܟod \���x�	A��ϡ�7D�6T�RE2^
 �rE}�+��9�>��<s{�z�;������}��0����=���*f"���ԓ���#~��	u����,��R��I�"n�G,��6�N���������ʝWt��t1~��Q�Jc|���#� |��#��?���K'���2V ������B7#�Y�����"(`�?�z
o�m����Q6<��u�mqD��-Œ��R�0�,heHQpS�4��G�$��b_b�(§�Z�D����I*���;��V�&�O��k����C��D?.z
��+mMf���ǃj��+M��z#�Qj�|x��52�?�J�W�#�Yg^g����0��d[�/�B��o�pf�Z ���:::�}�7��ȕ��&��14b�q�O�BT����j�S�J����Gã����c�m���_E���
��&�y�s����CqUg=>�zF�Lh�&3a�]d�%��h�As����⎷@O��Wz@�:��l��h�uw�ȭ6�M�&���+��.�uS�L�%�g�X���bL�y4����.ҏ��1`�VJOm�v0��g.k��'UY�����ۊv¿*�8���R����O�/x�J2���.�S���EB���$���Vky;b]{��pu�J�t��\<֧�z:�Q�K�=R�s��{B��$����jhO
�������A���ƫ��0�������B���qϗ2��f��c�+E{�#U`�Y������S�^v���D�،K8Ѹx8}M¢�����O{u޸���/��oCZ��vx�!_-wo�	�6!4��!�ՠc�����5ȥ��4��7ͨ���!4r�hUؕ�/�Fǅ�v.�ݴ�á��"c�7gX`��3Lǻ��k��O�z�)�̛�Z7PV7ny��UUA-�[d��!���	Ԅ�rшߘ���t�oBPý�x�n���ƊB,� c�]�y����R����Ζ���y���z�r�-J��T��/P��o��p�F����|wt:6	�����1L��|3?���6+�W�~֌U��;���D�y�^����Z�%"�?*�#z�ģ�
�VPi	���_����v��锂�kDO5_P�܅(*h]��*�,�V��a�2�>��=II"�Jm�}W��s��7��<V_�h�v����yq�NV�^9�]CN�e�LfT%���3�� 0`aPL�~�З {R��!��6���b*�M�z8�Xي�e�d��b��Y�v��OO�%c�;����a��RO �t��&����_olǡ��H��]4YC^��[<C��E_��Qb��Pl@����G`�R#�����Jk1$� �Vr'q��Ёs���bD���x�k_�:O����l4 ���m�.����7��&���K��3c4�	����ǫ����SIˇ�}��g�:�jݶ�г�ȅ��q.8H��a�r�e�`,b4�1�5*���[����n"WƴnO	�7��8裌4P�rS��`��yv� p�2mB�˙��b)����d]07�^}�ީ<�y���K����"��`�5���ԑ��nIMǕ7b���c&�&I��*~j�^Վt��}�d�t�N�\_*�����E��>�+A�������3YBJ^���,����鉶�R�Ҝ,T�&�(�T�tC��ŕ$DL?��ԕ���kyjߚodSW���H{�ESy:*���{]�)򾍄��D/-�P�5h������h�8��:璑����rM�n�c��k��s�@B(����P�\�\��T�)j)L���A�[��KQǟm�^��d�;e��\w}�o|.�V.(\�ĭ	fZ�uOPۿw�Y���e���j{f[���<U��E|%�і��Q�6χ� !�D�^/���=�e	�G�2��4�����F%#njq�y*��8��q���F��<?�pSW�����V1���n�וz9�rICУ�^��"aZ�:�1�wo���*����� ���H%�!�[2��S�LJ���X�lTc��uy�W��#����N�R��<���W�)������ꠚk���m��7|O���0uCc����l�H�ٌQ�C_^��;��4��Z|��d>�yK~��~N�N`��|&����`x�=B�?��4h��\K���x/g�kާՕ����Y6���*l��0S'x3�L�4�����	��!A<�Mr8��9h��1���#�]�ގ6w����Sl�B�	�2ֻ�
�ӂjXkla
�:Qy���F��F�:;QXup:|J�+U^�:0Rk`ɮ1�+�)�s�B�1R�}�rkT��3<V�]=�������O��I����L돻��$��Xc��)B�Q�h%�Lb�
Hۃ�x��V�O�c��(|*`��l7Xi�sh*��Z{.����
��p	�q,nł��!�K\Ŵh��CGR�m!N�]�Z��R��ֲz��?�+uGGi�<a�}��l5O���;���U��1Q��DR+�)�C|�O|�-F3-�I0�8�Z�%9�"�|�"�hhs{�КX�р�t_�]�x�{^�&EihQ�+6L�?(0Q�GOD��66�	B�΢Y����d��V�|Ae�� ᵦ��$3�S���b��5������i.瞥qU���-�?��<M�n��yE$4��8�;B�?T�1�����l�r��hE�*�ۆ�?U� �K�3�l�7���n�Q��z��6u�3�\WHwɪ��w��K"	Ve�Z�_���+�*��+�2O��.A�8K���*�\}�v\/$��z���_b���9�<&I2�����D�7z^�nͦ�#.��L(8m�|�d�����\ޘ�v�UL�j̥��Ҭ�:�,�'k�؏�M��ط�]؉�AU	�!�RK�ۣ���k�}<)M��*��!�����ذ��iڗ��̍V�i	��mJk���|��D0w#�]
�G��U'$�Kwp9vɉ}������!Vۙ�s�톿�B�����%��U�O�&sl�.񳴴��40�Ei��صG���caN�F���D��n(J2�6"$H̸ʇ�H�5��I~�0U~I<��!|��!S�x2:���m��`	��)]z��<U���`�#�-�iK�^�}KP���j����O%7k���sW��>p���pU
��⍼Y��6��o�]C�:8��M�~$Ɇ?_�:pw�����?�R�-c��m�ώ&	����n[Zp��bC�7�j[G	���Z�h4۟��M�8�<ܺ���ЃJ�L��Y�3HU�cR�o�+p�g`�5|���;>��Q�
`�<��yÿz�>��#_���q�!h��Շ=B0��s���(*@�gX;=�l��Pt� \ڠ?�@�mB�|ոS;��/�}mؐ��P���'`������p�Y�S1<v���9��VL���@���a��ً��r�M�{q;%�0vw�U�\w�r�RJ�E��DPg��(D���ʈ'���ơ�Sʢ���z�<_�e�nk�v����/��a�hZ����O�/�o��v}���+�k�3�P�)�Ժ>L����]
��GXl����J���#��m
��l�7_p�����d��r�|S��-	��j~j ;��
�{@@��?�-�'�`�����Bg����8t-��C8� ����43g����1dD�~���=f���-e��eq_2�W0�?����۲7��� �:��-+�։�+k}K^m|���B���l~�|��U���|:2,���l��mIwrM��2s�=�회�K��$b���Tu����説��_E}�w�P�<B��>�a��>�F��������v�*����>��v�pI]�[�����jZζ�?��Ӕ�}6o�� �� ��Ī�ko��S�����qy�`2xwqNY� %���h7�� (VmDzI���ӭ��us/l&��uL������؍P� SȆ��n�,����%9]���"�Ԥ�y��31�_�Z+f��y˘�c����] �]��=v
T��L��p��3���a�tk�H�6�Ò3+ڬ=Y�6Af~U�ᵷ��Bt��~z��H���'�. ,r��,�v�-����n��@~��0��%��
L���[O�k�y�p�U�TxR$�O��v8����W�s?S��H��{��k���*�͈�͖��t�nB���P�����@�T�
�(	h߭ޥ�V�b�@U�jjL;�;��_1 ��/�#m�J0�)4ʀ/d��#�S�	#����٪���Vg�*��+��w�G$�s���L���ݠ�缯��1n�'ܹ,Z$S9cv�
��A�eu:`����$fC��s���Hu,)���Qҵ�4�k��D!f�I��ӱ��{h��*��~֨��yi/�NJ9u~t)����^ŏ�w"�8�7oy^�2��׹$*J���MB��ɾ�ZY���~+5I[�TV�1h������1��F�?4OM2qZ�v>Ә��?�G���"�w�
�"6<�&��ꏉy��b�+o���H+Q��ɖ6���akQ�"`�$�.(K���o y���F�����Jm#̸&h2���Pp�ȽBꢼ^�o��C�_��^�$����.f��G:��V&�2E�OZS� �����+��z�h4���ul*c2朥��@L���}���=�Z�hB��J]PC�����7�ޜ�+�g�b�����d�V�F)ʹ����?Q�y%Z���3%}����X����ax�0>�}m�A��L��GyLGpTC�\�������jRIC�KaY��fɂ��qۓ�d�i��#N7)CA��%�YKo�{U�ߦD���0��}�ⱔ]E��@.\��p��%?as]�	�?7��*�q�|:ӡ֌��ir��@�B�$c�/������z&��"gU8Ŵ��/z�
�9B��vAE��̴�M�H~���ß��ae��� ��H�z1(�U����Րv����JX��SF	����pÇ�s3P���4r�&|U�x��]��;��0�DO�N��F�E��M���«-�#��qT��^�hp���C�7�K�(ں��0�O�߫�~�c*�ɯ��10���^��(��\&���q��>��d\��b�pc�JM	��QuGL鏿5���[��8B��=���8���w��i�y�4�^�zwbR��� ��O�_���6nT{/��?O͸!��v���@��A��c�,�8l�����`	��R6�8Օ�?n�Ͽc�Oߨ{���,�p�9�����<*�^���Vb���S�(�"��I|x�� ��3�H�`�������R���)t/<ՇKVD������^J]�iz]4� �#x��Uy��K�Q��j�
��\��NSRl	��z���Mÿ�ɤ�{��OU�_#S��4�$k.��S'�t%�kYeT��?��s���1,X��Rz&�{.aP���aS�0��Y���j�-��$�?W��Y��~~���n�$I �c��8�b�%�Fq�l/���1��}r$%���n�h�N��@t�?b���=�mp�x��y�^�6������{�E0������	�%�}��ß��g�DY�ͳ! �疋)�r�d���a*ՙ�@Ư�ư��~�陧9���}�O_�%N�9�OF�n���C����H:�2XLZV7���a��d��>Dr@����w�6ЬUz�����z�#�ȃ�p�Oj��A�-Js/+͓5u�9�?��ǫ�]���j���;��O�q`�'S��:ƙ������e��#f-ptddp��X}\v{8��ܤ��C�"���e�p��/�w� �[� ^���m�U�;+d=ESx��s?�h`h�i��	'�@����~���\>_�����{'L����r�}	�,bԬ���1���>fB<Q�����p�LdYm����״�c׽���A|��9�y<Qɡv�/���)�]f��o8�U�R�;v�i�r����qgq�3�Mv�/���2^��ѹ�p����=4
u}�(��qS|9���z���E�;D���$��5Β.w��&���5+ �^�n�w��U�S��'D���,C�fW�H��� fps��|h�}�k��J��/� �;���<"��oM��y=t�:��PP�V]�(�@�S�%\�vF@�o����t��{��z�Jk�LI�k?��撵n(��hΦdF��ٌ�4">BM����YӖ�Ll0���M}ZCB�qs{TCf���m�%s��q'ɺ;��Po+#-X�����Umj��Ca���hg�%�Z~djN��`�9�M��BK�[B������(��mu�.�����Z��Mi(P�� �xM�Y��Y���`sflА���K��KX�Z!ї��lQ�9;nxLH��s`����u��Ն5�K������P�$Mu���Y���ب�\������8}n]�	j�ެ����z'
��W�If��BF��*�����Ŏ�:N���5�&�9���߾�A��;m��d��W��O�3v.�-p�f�ι�d����2&�� ~u�{�ށ�0��$eh�taS"�����5�,ˣI�*�`���8Z�9���1�,��+����K�a��n���_��z��C[��(ĭ��K��� �g֗��,$]{�S�Ll��� �9Y�y�n��W1@��JP��K��"�#B%�S e��NBl_��˚��^�"�e�CĈ\� �t��'0;Ϝ��P�|��ǜ8k��3�b�ҥ�N�d�*(�*���Jj�|r�I���;"�; �)r�d#&ąx1�TW��x�ZfҒ��C�8'1��Vv��H��u�?[�W�,���+��' �j����J엪���{�1�R}��+�-�N�l���|��KgNOt#���f_]q����6L �U�WF������2b�쌤E�0�(�f*nB���U��!����[ r&A� �뒿�%�?f�HnM���.Y)��H$]���j����u[<��~�E�IaE���_E�&�Do�W�l"EW��kj�5�m4c���G�l�r��Cp�
W�`>�i�
8O�<$;��@��`�i�r)F9��9;�0��R������k�T m��mђ6�|�G	����n{�%+�Q��R,/~����|�e'��e"F�"���ͩ� /N(����ئ���ቧɷFN�q|>�]�Y�jG�_npO�ƒ�,�B�#�'7��H@���T�^?M�2,��L�α�`0mc���@�����j�]�!�xlJY%�{�hJW'�;E�.�dƅ��U�$锍T��U���ǡƷ_�ɀ�+��#v0�{�lRM���_��d��hj��X� i�? w��,s�������F�Y8�98yTP���"
$����I�ݐ�T���W��9w;�p]�R��Reŉ�ȧ�$p�u����j�Ͼ���	�^���,7�,��N��7n=t�>��C��|��UcI�\�Yքc: e�%n�������
`?t�����j��@&�w@����Ɖ�c��yn�׻�	�'���>V'��� K���X}�/L�0:GϳDO�S�8���Q�\Ѝ'�����0J��Rؑ��&D8m:2��;@N<�a:�%C�^n���[:M����:]9Ҏ���D�gsJ�Ԃ���ӛ���9��[_��Y�|���"�g��%_^Ƕ����?`��<�M�s���Wb6��.�f���ġ�����ˈ��=��숩̿�G�3GW�ö�t��Hr����UH�"��������08��+������`�I��Ǳ�)V��@x���o�qu�%�?��P+F�U���X�P�{Q7���I��@��ۑ�^_G��XL���n.��MPK��"�7X�uRx�SA��D���zY/k*�DH��N�(W�R������X�q��a��}k#eK�j~@�����F��M��6<=� �V�\Ov4���ʤr��N_D�!�㼘�����@���r��&�O�����,�1�B0��itC�'4ޡJk,)wC���0?��-O
���x�qQ�W�n�Ԏ���~%O}	��1�=��mu�ӑwE�0�j�0UO� �����e=�hG��%���i�8����h���cڀM
6�Hκj�RPI~jz����W<��v1qT���`!�����>��R���I�k��o�m�w(��?�rk��K[���|~���/)�w�R=�����e����Y�Ŵ�i�d����fv��?J{�1<`s��$"�@Q� ��z�&_�?� fQ�u8i�'��8#X��c��SCU��d��ÚG�����jz��ט��Z�-n:x����qMZ��]�>����+Nج�Z��Q@������V��
{�_a
R�z�JS�w܀%l~T���@�R���*���.�E �^1�F�J7"�V�'����
O�A�2���ь2�JaБ1��jpX���r/C��&���t�k�I�	�}��d���B��t�m^��d�c�%�$P��9�Rŕ�3F�g�-Y9�̲j�t�	"�̱����tλ����!��Ą@�^Z�/_�������b˸��sZ��7�O��z���j��k�3D��x�8�2'���|��-p�&s����Y��䙼{}%{��my�D����w�GL �OC�bM��y�F�)$��HbT�^�M��
�"'��`7���bdG�����R#R�DW)X1���Y�,dR�r\�Q"hE�T���xnd�0(z�4�m���e�I�����o��%�'�~��>M7�7ibXR���A������)h��!�o�bXz�vay�=E��,��ς�Ď]iSܣ6.���]:��v�[C��.}���ۃD�z�n	n�[���܉�%�VF���]���jW��D��8���d�n�d��%�a`M�;�'��Vv��]�F���Gr� "b���&���:61e���bJ��1�_BT��}ĳ�|��
���[no,�Dx?��[��U	����9�3Y�QUi%�8��2QB�?��	s�~�b2ۤJ�t-�կ��EL�:�HM1�� e�Ӻ�ӱ����$+����'�a��4�d�7��<uc�3IFq�d���y�9s��0��~\�s!k1�(��:5���_�R>���zVrfeWY�d�C��}ߔ�fv��Jno����0e�>����9*������s�1CN\+��1�KJA�i�,d���?]�)�9t7�,=a �V	��	/w���T(ba��l<�x^���l@��@Y\ҙ^y5%��~���/�����\�\��:/�W�����3r�mc�X}�H�����_��?J�����	ގ
�e���A8x�l%d�o��0#�&��j�}�j����V�9:F bU�E���M]��nx�j�����5���3cihγ�;y���I�_	�O�$m+�x׹�{�2�$�ͬ>xI!^���9��(����ݝ��$~>��	���xP��d;;MՀ1�ԘS���X���Ew���6���0�����e3okldЧZ<���r�2��}�gA:=K՞1����t��ȥ�/��DV�/_���>�8W[���\�G��"�����-� �;re�6>L׈{/1����y�Q��8 B�-�8ٕ�Lߩ?��p�}�`Z d5��`�8����U{
]��ᯆ�eh�r��gXVC�"�-�ՙ������A��C����|�(R�������)8Zu������]u�����3+q窴|�0�ѯF���;��b�Z��O0�<�o9�5"w��HI�rmR��m�S�[�A��jw#B���9����7��{eeS��˓Ϙط@ =|e����ڮ�<ܯ��cu7��	<�k�3:̟��o��痔`+�@�G�c��2:qm����z֬�`��/f�	���X����/c��ڊ�N�Z.�I�7=N�"]��k�H�(�f۶���#2�B�1�w�c�ث���lp}6on{}6���d�ɜv!(�g�񍪕�^�k0{�+�����ٔ��̬T�W��[F�2��>"
��J�k� [�nG�������T���(�<�����dѕ���&z��_z6��Lp"G��e�೿� ,�.�e̳� �Wt��,8��l}�nNW��=���P0�:E���"I?Nn���pi��$V�D�\C�_�}��qp����,�g,���I".�/�T�'���jƜ�`Y͸)_b��h����%.�R��F/T����,!�[]�l��'_0����l$�Ю�K�j##_p<��W}n)֌���D�$+�0����<�N���X�_q�2U��ʛ�i�i oxyڎ�^�)��4�Wb�װ���E���;O2SrY��-~��Y�[�Op$���B�Y��Mjg��Q�Bcs�W�ϛ|C�5����"�"��	j�*g�~ �1��Mɲ�ql?�������d�t�a8s!��2'��n��7�U0znF|m�X����2U����]�����[z�N��[Mitg��
i��w����Tw�����h�����􇪑$���(��@)':F������y�:���3�ڥ����+z����{�b~� ����6�x���]P��J�X*Q�W�K��q���g�ȗ3)~���p��W�9�(7��A�!*��;�L���[��+s1�P:��z��1�NP�G,������p���\��.��蠈��i.`���yT˞���4�jd�d)�G�
)<��S����OY��H�\���y�&��0;��f���K*6H�Oۡ�r%��=#��A�r@�H���%�adI��K�%�c,�U�� }S�6�,����o��I�S-�{���)�{�f]4"Ű�Apm���W�7��¥�4�m�����q[�[��#���f�[��*D�&yO��2!Jq̇wEZ-75:xƶɦ��y��n��u?���!%�	�F��9�H�i��ޕ�k����<Oi�1Tk���l���ƹ0%U�]L�aKz^3�8:3d�b��64S'Hp���rV���� md�f����NdU��}�0��{oE���yN���4>����*�5PH+�����6���P-�g����U8q�g��@�?��vm-L3;��#^�X|�C\�g�£�ӂX�KK�,{+�v�f����Y��"mL�����BKJ�M�s�/�LL5���Y�ס���q�Ó�M�
V��������mW����^P��r�R�]���/@�=Z&��C�]D�D��?�]`��Jr��ž��R�Tl��3w�\K�^�8���-*Z�b�uv=��c����;o����o�!2z�v[$��Z��q24�0=�V�쮜��`4�Y��j�Y���>ɲ��0]+0,C�Sg+���9ș5�\��y������G��*{��9#�o$�`)pO�tJ��ې��O��(�xhb�8�h�v�9���Qrw������1��m��i.�0����R�`��Dm�_'�@	�{��=0Eꓓ��T�+�H��6G1r�B��H���c_n�mc�ښ��D����?�Nh�|&{�+��8$1&G=�4���3���>�Tڏ=�#~:+�����H�S�����,�rd�G����&�PM�6��(tO�w[-0�v��_P���֜�a�|�bbR*evT�X=�<�w�(�:�ih�b���E����a�T$f<�'���3� C�����T���@�&�H���I��i���52c��kW/���g��^�����������gc�Q��KBh����Q�U-T必Q���"�[.�NgqbH�4� ���i�\O����g� h�r�ړ���~
� �C{�}��^G3������:���1fb��kE�J.?��������j]V�I��2'~z�μi�)P��V�\�Rֈ<LlM�%�U؅�����4�!�HV̞�&������XD�<M�ke`|�d���!�>�]� {��޾b����!/�� �����l������KΕո��z�[�^���L){I�oe�7Na�E��ȗcyVC����[������f�������
�{�2YԴ��ґ3lU�p��H�Nt�,��/n-�'NS)d� 'j9�(򏈢��ы���0#��ӏ����R���{�ڡ�1݉z]�����oo?��K�G`��;��[
J���K�����ܿ������)�K:�]]�&��!+*�R2-g\���&إ9��vh��h(�|�����_�V��z �eY[ ��d��?���U��i]ŗ�1{lvy^~Nh4L���+����r~)ğ�Qra�9) �,��������K��f|������@�D/`)��:�y���^��(��,���2��'^�}�&�+.��6�<��O��c��?	 �ot�����-���+�����;S}fB@��Zy�k�w-S��\�����[��l�8"?2n:ٕ�E��sP�btű�(@x���y��<�!9�6�$3 �Y����g8���%��;�w4����Y�%	kT���m��r5p��J��ׄ�`����"jw#K����p Bf�荢ZV�����.�̡ ��S|��d�!�VEz�K>k��`w�������v}[8,=��T;��M�:70t}�
u�ӏ� g�l���r����Oqt��R��m�X&��!�"]8Y��(�����H=7�
��Xo�D�g�����f1C��+��T�-X�&�ֱ�c�MCs|���_�}��)oT�/���D��8Ń#���_�J1���Ԃ�ˣ�+�������p���f=��ٿ�)B~������M��m-[�*}�^�6 ��6SiK�P�����-X�9'����$
o�����,�O�SG}	P�S�>� �M�ͫ�~�lmL�9���,�9p��K7h�=p���9q��2�(���	�~������-S
�n��ZQD�r;�A�Zz�m�U��@9Ϩ������|/�����*7�FxM�E�k��5
#ͼs�.Oʌ�#v�A����FM1�ܮ��a�nMv�����l��ƾ1�������� �x�NRz`������w3ن�ƅ���A��Y�?{�/��L/݋}tn��Zw絚�껠���=8ۣh}Եg��x�ziydyu��iۅ��-svD�Q*��F���>�����������v��P���8���UT�a�z{�9m��߾rĤ��G�����a��cfHd��j*+.49W���e��V�+����Q292t�Y�M�JB����VB*ᒬ<�0���(l@��NWy}�ɻ��X�nM˟��o��M�uE��廓-��j8���;��n�����_'�SMգ������F�Kױ����3���`��J"��0Q&���)*���`��oC&#NQ͢���%�h�����!�,8���Ê�؎P�⟇�Ij����_wF���s6%�Zk�֞���P�1c�\�C�&�e;'-����-�,�`�����YXp�z2=H���l#����:���S�c侳�q��ƙ���ٱ`0����K�LX�U9�?�q�>�:�5�����݇�U��S�|�I}Σ�����q6�8�R��(��f�U�<�E��@£D���U@J�i ��pT`s�2�^�]�2b�rO��̶�!\�~i��[qF��ob��?z6Q3([���T~�n�2��>ğ� &��8RWޞ��iW�p��#��[��?��nM���˫�H�� �Y�̀Fɢ/�����	v8{��V�o���N9x�N��V�ƄM�v����-�4;���Dq� �ޤ�HByT�{`S��+�����j��NJWM���<6}̒{��$h�ߚ�;��8��>�,;�������LJ����q#�y��;���5�8��p�L�E����.8xΉl�}�9jV|�c��z��*��%�V���mK#��h��:���6�%j��(a[�6�������ovq�]����9���~>���Vڴ���Q½=ɛՈ�ɐ��"#�&2�^��be��]#,j{���v".%���EW1�����b�^+�@c��D��u=��3��I�b`��"#9F�������F ���*�S�a�,����:�� ���	<5H��]�+,�����i8�#yX�S<)<k��{f��G�/n�����,M@�	_�u�o[�����##2א�)�K[(Ӎ�p�o�ӟ0rȔd�6����4���\ɠ���Q9�28�H	؏u>�/��4��	��J��e��ʁ�0W�}�0�?�y���8	gw�%co|���O1g��0w��|^0�'��)ln�}�W||,��̵��s���q�%�o^q��[)�wW��iyK&�J�;D�W!#�kg�*��9�x�����'�1UpT
��\�kA��(N6;��]�.��|qr��d[��h��h�Lb/�����.�a$��K��zH �E�d8>Qy�wis���Ѿ���S����B=�(3C �$*Pv��8e�+H]�&">��Tݬ[��0�@�a��?�mE�)t�K�f��!�s'Y�C�tw�}yQ6۝����og[���U�� "|Fq|��L�9��q:3T�k?��Ӱ[F�'�zw�Z�9"I{(%1} �wэ<}�k����C�����Ǔ.nS��-��	���/'3�t�Z��!�Z�2���[�����>z�H�	D���7ǽ `W�P�q�Q	�|�\��<_�`��3huǩ9�:rr�bZA�S�D͖��gۜ��-枹fի�N�q �Ɛ�;$1I����6��[�S.���G�[:_���jN�������4���҇���l�Bt���LT��|FZz*	ږ�5W����#%n`�C\JK�����|`�F��^`\�s%�㧇�[O�k�s����4�Q
'm��+��$s�g%�ty� ω�̊I��期5m$���@��3xd<�/	����Ͻ$`M�!ى���n����A5Hk� b'gIq?6$�
6��/ؾ&px�ӵ�3�#�g��p�4��g��"���C���Ĭ�c�����V
���WhL�Ҥ�Yx��#��t�7a����\{��ҝ�ڊ�E�rsL"�o)*��v�H�m�cI��@�->��0ۇ��/ʏ����)���x�qdwAO��?��������d"2�m.\�w?����{
C7�es��H3�粯���~~�LpF#�n��)��e�>�T�`�鯳Ԟ>D��z�D�����~���Cs��mO'|����o<�ߨ�G)�*��U��$r#���bl$K3�Pv�uH������ț���
^��y�6��e< w�Ԯ���)��z�ZVN.:����V�42�3�o�5g�$��u�����(���PU&��+�{�i�k�� �қ��ʀ��M*�����Xyn��$��V�K.9Bp�0�u�����ػRf*^�K���4�3<KV�G1��I��m��i�s���;�52m�-Q�0�!OwEme�����K-N��ԕ��.�@?{wL�+h�nbq�"$1+0�\��tG��c��p�q�-jT<�19r�M4s�i��?yY�������R.��+b��i�x�Cx��p��c�Ő�g����y��P)��b�N�-�$��X�m��+��@_�ew�w�
;��]�\��0�om/��`ȝ�V�Hw��n���5��u�!w0<�S��:�y�>(+�2�U �sl�O����ى�� ���@i����m
�~�P��3,~C��h<�������JX�inm�v�"z9
Qf��ɼ0��E��b��[!��p];i�g�Ǵ�Q�\;�E�,�7�E/N��ݶ��C .���@���&tx�}['��}�=��c�^�$�ͅ�|�i9�-B[j�E�Μ(FrN���N׫�0�4�-{;�Wqs����M��4��L6&8�㺓����_�9 pYE�;y�0�N��xK�\�&�~φu�hr÷&�a������ם'�Kp��P�ƽ�qAʲ���G��hD4?�^9�[9��!VԞ��G�2����&�=-9\�XO�S8=&(����z�Սa*��q&��E��Y$�@��#!2Ӏ�N��r��a(����rG�WP�俞�!����>�X	�� ���Xb��f9F!3J��w��e-���[��*�->Y�%���<�#_�W+�$[�m�p�%�_z�FF���.f�X+��X��d|�Q��A���V�m,���*�&':7ϗ#�&�VwF���$q�,�4��5�����!��'�y;D�� B��>kS�^�)t\�b�U���cNUҊ��`&�@_��B��R����4Cn���ĥ�2��9+Ѵ�����B�N��̐l"q�k]�	��e^.�X��d9��7$�]�q9���.�A�� ��z��%�8��#���kM�J*$�
R�+�����iF�����_��*�g��� {C!��d���3�o|b��t�% �2=�Rt<)x9i-/���F����Z��H;yD7.&�CV���t�!����fzh�\e�1j��j��_�`�Bo�Fp�}?��2���Q�\3�^?���a'H�Ns�翗9c�]�D/�͆gM�~�g���U)Z����% h����QNiC��.c��t�0!U�E+p��hK[i�"'D��a�瀍�XO�۞7z1��ؠr�i�oI*�k�J%�h§r;��H< [X�,���m�;5?{VfV�Ҳ��;[���Lia^���#�J�_h�ޘ���-�RY6wM�&0��?�}��jx���"�_� �^�V`��/�e�Z��g�`-��� ��	?OR�8�~���~��!�41,kiA?�"�x�{-���I��|��KA�g�Wg��z����CӃm*`>����n�x��*��~M�g��#}��������eEO4
U����JN����,n�^&'5���X#"�d�����\�L�/��~A�&�x���q�c�QL��F�J��m��LV�ћk��Iq�S���)� K~+�%���G(6"� ظ�7%��w$���
���d5�9!����))�|��C?�ˉqN,���wi���ȟ���lEcHz��n�i��#�$��38�4�|���3�
��'� q}���I:��b�]A���ʠ�7�Ɓ�|7��.�Q��:��d���[i�Vw$��Ć�Z#��sj���qW��bj��g!d��#��`�RH�]�B4����dH|�,�[���I��|�k=s��i;�v;�O3���T{����C��B���&�P�c���*
\	D��ԃ����rp��a��M�����O�`��+"��Hl���kmu�����6{<�o���gC�P�d_���	X��*����ơb�5H�qC4�j��1>����#yI�h�9D{�G���Ǧ.�*�"��U�i{���yJ�.�W"P-ZB���v\�v�!_�/�ʉ/_Qĝ��`��ڰ2#̪��D�b{9ӆ������l�GKi�j�|WT��(�Q_�6������^SP�dCu�T�@ŧ7zQ���2�~đ;S��u�2��Ŕ�]��p���2�}u�K�¶8Sʹ�A�;��T	�b�,*���;�=�,�)�:=OH�LW�إ�lXz��+�k,%�HU�';},�/���R�����=�'o �hb�ab����8Q��MWX2��q r�s��\�68�Ĭ�\Y>\�dEp>ZJβ�%h,f�Kz�K��Ե�6�Hn�a��1�s�3�M�a���QGř[�P�^(��+��؉�����r缫�N������dk�V�~cP������F���X�A�n�Z[j�J���'nJ�+2~�ΎM�{�J[�Oh����LS�p<H�a������Z]�����JK]� �ݸ�>�������	!}�	�{�`��&IK)���Ǔ!�۶�6ZILp|��W�Z������a��ϐL�y��!���9�8�0��sfbw*��	����u�X��rm��Ĥ�vT�R6���Ȅ�7��U�g
�r�m|�[�?Q}�ٙ�Ҽ�ݎ:̿p��]2B�(��3�����$g���!�lA��Ka�鲯�C,> wJ��R�$�U2�~DW�x�=R�|���L �־���7�M��sT����oT]�6y�?�������H���U78Ox��/�V��໶f/���	�~�	kq�E���u��J�$����eL��\�g�t��=�H�]_@����-n����9U>�΢�c}�%��:1(Pw���έیT�K���h{��^��]��v���C��[���?�����H�?�cE	tp:�*��e��h��������ƍe��?��'c�+�f��0~�;��`�S��9W�oNU�M��؎9�:�V�=eN���s�������s�Ӗ+,rZkǻ���_))W����%�
@�G����g\K(�,W7s�	)^��xI��tV�>��d�1���7h%ߌeEt<�G�;�V�݊����}��Ι���n�V��He�o�?�D:��Ȓ���tCq�o�*&�f7{�ƟjBj\��6i��qec�,���y�����4�v#�>HU�@E��&K|�)�o�� �!�IL #�-�~����V�b���P[��)������i6:�����7�F�/ƐH�4֛(VL�i�r$I3]��������8�@ V<n�r��vr�Թ�l��2��bb�v�G�!T�D|̥�AB�4E�4�~a�^��Y�����e#��؏��7WD1K~��!���qr���T��A-����Ԉ
�!�p�ʩ���}���{���5��(�p(^ ���2v^��<��'��$�9�Σ��.���v����N�' ߶�5 ���^ k�W�O�6��@�O>g]��a��ݚ����<2���\�TR���m#�)(b|֝�7m���פ텭3�wKZG�V��$j �}�eK��Z}e]�x��-��=x�;��.:����L�ߖ�r����-7�mnG�Qm�:�j7 �qT�cz�ت��PԠ]�j�ci����h�k��}��ތ���Gu
�P��fZ@I\��Y�e���y��$�#�-Sd���Y�����m<�+]gY�)��e�]�!��3�ǚ�{B�Ҟ hA��Rp��
e0��ARZ(��\I��@�Y'5�?54r�b��=��z�;�!�O�'�����1f�)FSƏ�;Ua�������G	5���2�u����ǰ(p��+�-��ό<۟UˢZ���o&p�S2���e�O�8p�"\�6ƌ��T��� ��1}Fz��y�m���x�R��⅕��D��Vm��'l�q��^��̏	H�V��|0f�St�5o�`� +O�"J�ފy����j�n1�L)#�e#��ߑ��[��b�F�W��x;<�z�?�I�8�s�.�y�'6��f���3���~�	J�J�$�2䰖�-��uF�pyS��,�-��R�P��Ik���	�m���?�[Ҷdu���F<�ь�� _uK��rk�.���Q�8ey����	(+��(kE��jEI�LT2�diARY4֞LC[�Bۉ#i ]�H^�)� �*]���|��YZ�L�#D��T�>51�i����4D^��43�;W���=��f��q,ydf�Okebo��`O���&ly�]���R�?�������Ȁ6��J�\�4�䝞��t�"Fbh��$+��*��N�	W|YA�X��TM�(Cm�A�]-�.�;�	��s�w�'��/an����AAq7�Y.[11  ��^!��bw�,`,���i��Ϩ��}}�����fh��Ջ����r�2>�ʒ�D��@c��@b���q��sF5�SFET����X��������}�tRhq�*� ��1��k�?Ѡ��]�����]qkw��׻�e�z�カ	;MD��գ�Ht4�@��ljx`���kX��v^�9����G�aCN��4�͸9���G)%h���3��� ��=��I��Q��ĢnM���\����7q���S A�)it���om�}�C�xV0�R�`Z� sɣ�Sf�nҗ�M����iê�	qH���(��a���%|Ǌ�����H�ۼ0��D������a~8ܖ,��mi����n;�3x&(�pf��	?����;��y�Ji���]��1�8/��6�����Cc��r�����t�DL�� �J`��a̦Hd7�]k=����ض�����_)�Wf[(��k:q��\�z�'��\�o��!Q���vż~yu�������q\mP.v�ao���2��*��?�bG�!������<	d�<�=��'-˄n=3H�u��uO���9�^����DQ��z��AƈK+
�Y?H�VW�;ހe9��<�nys�/�cb#���#�����e͸c{4FQ�-6�QB�<��#�`�mX��z��8}m�gN{�fL*8�3�;T+�����>�)y卢�2L���-��a���)��CKYI��J�?D@��/�}�� �`�Y0���ȳ����#��Z�9�k��a�5\�3�t�ii���1�v����4�-7?Ĉ��h�d�8���dB'�N�Z�u����g���L���D�̴Aq���������[Rn{m���?������L�=W�m<�|�b���?|0�-���Q�ĄK����DHu?�DU9�|T�Oh��{�Dh�Quʺ�O�eVT��^p� 룤4J\���w�Zk��`�XD3�ʛ�`��g�gf=����2l�_�T��,w�kFv"բ ���bDd]Q_��h+^#��w&��K�������֛v͇�8�[�)r׹��ciTH�ڌ�'{do�U��dǭIf��O��M�����b��tB󀨑���G!k9�Er��a�=��y{:Ů� ?����68Eacـ2��7��-Kn P$t���]��a�I�l�Md��qs��n���D�l�����/^�g�o�â�Z�miҜ��0\��.���#�}�b�j�J��$۱b,��0W��;��N�+^1�y��aR���f�H��v�W��57��* ��S%%��R^qRwu<M<�%�-%�R�S{�lؚ��J��un���Xf ��P;����	O8�����Ӏ��D��&�zm���H�+JP���bmo���)���O�|����k����ޫ��ͱ�����T���������H��Z�7A���#t���UN�FB���Ş�P_rgй�D � �E�|�:`�t���?r�J������hD�K��{T�k+��{гVh��'6�>�XY����櫥��f����
u�fb�~�de�m�̀V�Bt����M-����Ֆ��Y�n\\a�٭�|��{si������i����t_2��D!a�ǂ��$o���k̿e�dF%�������e�����:�����	'sW���1�����/����	���BGI�~e	A�4�^�P|�_Y@�q�r��J(��B�F,-���}b�I��sw���T��WK�I���N���M�v\-jӰ��c����cp|�{T��ܱ���a�qY�ȷjFS��z5��FU�G��Ye�����4�z���qT�ФP�hR})�:�e�������ʡ�9[-�x,7�s�M"G���\���V�,32����n6����w:
��l�
H�7�8���n��NdH�l�<�]��6J���dwv˨`��V���m�w���N���5�։5:�?ʽ� �mP,��3~�q�X�WDc�xQJ#�0��-�u�:�֠�7'��͑��T���W}���m���~$��.����	p{�S� �-��t����������� �GR�p4�����a�<���/��?�N�w�5sl�O��i�п������_~�m?*���s�4PHlk͝�-����HLV�
h�A���=
>�ovc����]l��VK��n�t���#�=�6����6r��t��_�21^��C�Uv��8���I�*� ��A?y�=�ˮpR#�➑�8V	�R�m�A��p�Kv)��`�D��i��?���<��F�4u`��k��r.)'�V&��`ئ�6�E�;�Q%��3ז�����M�����bA$0���[`=�B��?9�%cIO ���0nhz�B�Y�L��d���A>���$��qLr( Ћ38ʨ��<C�Q����1���9d0=�c@�-���s�Q�g/�!��j����\�dh(�:�gt��8oC�5������,�\�����ռ�8J�[�����L��(+q����$ts��|��0��׍J�:�Xw����skK|-T[.��A���D�g�Q���ʢ&���P�""� 󏺡C�}} WKM"���> �j@ Cr^h#M-�m�Œ�Z̵lꙞ��:�+��[i���.4~z��`1��`��>����&B� -%g�+`z���_AƮ���%�����Bu
���r3��	�%3��S��2��/Pk%w�K��i��ó5n�оа�,q�&r���y����}�LQ}����slR�γJ!
tW�t2�ͪ�$qJ�1�پ�����/NV��H48�	�ת��	��^�dX�����h�Sv���G}�;)ʕ��������@�A>Nm�R�ɊJ
۹f�W��*�+m|ԫP�ɣy����Nq���d�v�7������<�Cy�$g���C�����0��>̗D�B�s���,RBg�g��С5��Ϟ9�z��v2�����9��`1A0��^c�����tp�QRR���6�4�(�iN��
{>(�f��d->��G�0�zV���<��G�M��Y�����1�kz�y%&]�V�����
e	cYt�7��\4"�_sN�yo�^6�o����6����K4�Y;�� l�d|�0C����f��Hr�8Y�7�5���Z���x���b�U�یbk�50К�q��H=�7|����x	�c�5Llb�uC;li��K|�\�[%a}�J��6;Yu0��w-]�T|m�j��Ǣ��_^�>O�B��@��_iw4���B��� ��\�h<@O�q�7i$��Y���ڐu^�7�8�RM�_n��?�y��4��!��#�팉={�(�ޅ��+�*��O�Q�m:%���opN�zj4�c�ĉ��vN72��fG\���!G�F�Nu���X�f�\Zؑ�x���b��J���.8�»����T4kY�S����qlSw��С'C~Z����&�Z�����F�'����
w�#��|� �o	��������]Ouz�ȍ��Km������F�b�����
J�����n\�&��M(q#�JP�B/0���Chy� ���<�{��h��e���L'�5��q�~�,<y!�83������G ct{
*x��h���Â��&ڭ����n��rZr���n|��'��2A�<��a�����g�n b����fhT8B�7 hcB�u�l��Hٹ�d��0S�,1/�L[dU҅�qV����xY�����fP��;����_��i.[D����D��\t�U;��������{J�t��{qQ�a8:�e����v2c�m&Rz��}�U\i;}�h��q��@���~߷HQh>�ӎ~=���𼶝������)�|�����-bƭ��^��+�k��7*u�2���3�	J.C��&4�0�O�t�64��Ű"��kIM�c��ڇvQ�I�1��ܙܷJw�-�� lg�!�T�@�<�Cl�XG�z�{{�'x��	0���l %�ZI�!X���;M�D�-�h�o�z���/dq�D?��u���ԙ�Dqi��aG�D�������y>w�`��όԗD��qt@���
`|�)��\�Us �CYE���hb�0?ؙ̗S%q�,������������#~�t��VY�)#!��xu�DB}�-�U�A�Rt�vxDO#9�>(`�c�w�ػ` ��ߨ�n��b��JoF�h�m6�&ש� 0�`x/z�8i9t��Ӌ��)�w��/V`	�
�naRxw�.Vtm�Y��Ԩɍ����Y�E}TB���A
>�23k�SU�@K�!f���Q'��X����V�\5��8����Q������#�$�\Z��z��h����`�_������q���ai�%8;��ڦ0o�W�qt�[�3Ĩ�R�6By���S���Z��?�Yܘ�Bі(�^����(�M+)ƅ�_�$������u�h�!�7-��l_U�?�^�G�K�d��0�?Bڶ�g���c2���d䉱8�P\#�2����!�hG���(�\��|�3T'(�l���1�-���q�  ��h�Wn�v��lM��C>RW�*�O�����4Ի$p��R��J��/�WFh_i�Z�J�"���=��OZX�>�d?��H�=�kƚd���#�4�hB�};a� �W��|��u��	���[�����,��X�ak�n|-[�� ��N?��x>�خ�e3�^�nV��%�$i��M��N�#W�*<���
���	���K���@_)���V�@$&�=\.˫@�����[i��J��{m��sg�)�/DC�օ���*���t/G��)=ߢ�]�`{҃�S��!�3E"<��l:Q���Iן�y��5u�Nkj؄x�g
I� ��г䲸y'(e�gW �.@��#��{�)+��vؤzf�6K��~-��ꆓ7E�wiK�T駮y���m9`�ɍ:,���+�-�j��`"�8�.�]��3ۢ�j�+��,x\�x��
L4�FE��̮�HS�(7��X\a�ѻ=�����$�>��G�u���P�4�D�5rt��2�8�?�@JR��>����p[Zl�&��Gq}�r8>W3*���
�tt�0����b^�W�ln�aߊ�U��آ��*R+���$�R�릳�}�X�DÝ��ߞ�1���"WM㌃7`�@1"�<���0�)j�'f�� �����f<�/\ǈ��F="
@ȏBK�K�'-P�%t0��+�a�l�
����=� ��\����_��Uq֚���Զ�t@./y?�D��(�-?/��,|K�C��C ���`����>̭̣P�y����R���gU>^���Y����6Q׹��L�u++e�x_��>�T����ҿ�O��q�'��	�^�����Y���@1xֹ�5>��\!ۏu�]�����7���0��^�5��;dD�]�C�%uя{.����~�8>��k�hk�{k+l^xo�a��Q~�A���J8h`?��w��?5��A������h*B�����'a��J&���g��5{ �ݟP: �6ߎ`J����8o�ݱ��K�vJ���[�P/lx�B2%��Z �8�I�yi䝵I׎�������3vH �n=`#y��#*�u��n�PUp����%��
�7�ެcJ6R�Ձ��D�,Z��c�T�,����G�z�!�ɜ���]2>K�=M�,�+(/1-���j��*H��H���
 ������%xq�4]��[�L�L�E�y��6=�oNz����ʸ�M��z�dA� ������xRT&�E/�<�';�Xt��â��4B���'�ڄ�Y��.�)Ġ�!CPN1���/Knu���2d�������+d�G�G��a�D��H��<̘��"�]ݪ-�9\��Ӑf�a
��sC��}�_.�8�͔�9�U� )�Zr���T��]
h��vÐ�ŤL�6�.!{�5;Rr"�T|�T�Z��Q�]U��e�}M�A�C� ve��]��X�i�y��b~��P��Y�vsR�y�O�n���U��ů �kԤ�V���� ;Q�s�:�ͺd}��7������z,6M�����"jC2���.�	���ȔTT�VY�Թ���~�Ӹ��;�*C����I�b�:���Sm�e|l��?�y��r��@�>o�����D�G�<O*�[0�o�����v|k�#�H�uz��pT���w<����#¢�t�/Y9�f��I�E?�ˑ2O�7���u%id�Y�k4���:��n�{���JoD5���c�UzO�j��h�C�4#�~��J[�w��&�J�o�Q��[.Dۻ�����l�bV�dݒ?��2)��0O�)>�g��j��?d���dn�(!ʱ�3�E�J��˰&a!��b<q]��AB2 ���R!�E�>��꜃�y��h����kG�w��`��a��g)��"D���jv��-|��g�2}�o26��.g�j�N�f[R���},���b0hѐH\��6��W��F���[e}ߺ軽�YDR�)��1P����"rh훦�6@{?;��X�P-K:� �*g� �|Qyݙ	�&��¨9F1=C2���w��V4ƍ,8��k����8dky���xJ�ě��p��.�ްҢ!=��yJ:n+h��EH4�\/ ��0Q[1�dQ�cп�:j��%J��es��mW���~���y0�d��n��Of�|�ʚn����u�\�{ݯ� ��/��{�^�j;�1Æ��{E�eJ�M�ZUw�*J_{W�M��e����~μ��#�%��CR�Oc5M2c��������1W��ʼ�]=ꈩg1
5�5�f��9�er_�SLB#І�.
�&}B�Z���w�`GC���J'�t�I���d�K�pg�6K�!i���WL��N���N~�"���W����H�&��_.�-E���ڄ�]�[�2�}�4>������c�t�t��j��˓T[o��VT��%雘��W4������nEc�A�n,��G����`h�G���x�^���0fv�O�,j�g{�A���_6��7�d������Ѷ�~��q	���=Y|,�^5����֟�N��(W|Y�ѳ��9y�3?�r�G7ƛԋU3	pl��N�U)���o*�(��`�
�۷Ue(5���G�ާ��V�a�F�}�����Rf�@�A��)ƃA��%��$},�V�ʸ�/��v���?�w�X�+��=Y�Jԁ��>�V3i"��9W���~��"DT�F��aZ�%�@���Lm�ˎ^�i��Դp�p��Lb$+ʋ;K�ѿi
5���K�Ga��Rw}n��f���6]���MFs��f�4�����3��������@+�{,b*pv�l�F��
��;��h��t�����V����`��`��;���7[��G�wMA� K���h�TE(�o�<���Q�e��p4|<�q��&l�3�g]�Bm>]�h���Cj�D?#�*)��{�,�sc*P�h�E�W��c��Cr�h�#���0Xu�o�
vu���%�l�`P6w������(' �P��s+��J��;2u=��"�����U�"�[�t�R�O�"�3�P�a���@m��X �9�l|11z�ϼ��N���Ǵs�{+V���a��?U��A�ޚ���襭s�VPĺ��!�)�גuX��`��Nv U�ߵA^����nU�O��s��Q]Z�i��)D 9�@��[�ay!�k��ɾ"��,�2�{�ǈr�N�<�v��.$حy��C�:�;/��AMV���%�q��k�&YZq���M�~�L�Y+��,� >nQ82����it�!�u�]t'DVE���6����^`ov̜���e=;��KH����n��1@�!�)�)*���M�c�2���#F൅> ��%���ذ���e��ؽ� �Xz� �{L!�N��3ɱ�]C�n�=�ݤ
ߙMʋ38�	�`Ւ%ۦ�)���bS1���V�<D��U���Yd��豊���W�i���got��b.hb_�
�(#�+��9��"fjX+�qҪW��u@�S�����H6?���{��6gS�=�-f��Mk�{�[2B������8k��,�T~Nh���Hr���k��×�a�BZ	d��;<�E�U*a�a�����j�QL�/2���-a�8�m9w�5(@F�����i���{���Y�T�5�-4������Cb�G�意|ŽMf�Ӣ������ k�����B����[�`(s/�$�!���C����������&�G˟f�Y�$c�<h �� 舳agee���?G����9�t�1�U�iXm'p���␙�4i��`z��M~�,!��g��$J�ߜ똹�5���ʪ�!yʮ-�m��VP�%����f�输�f5֤�E�r���	l��+�&�o"�!��"�x�ó0R�
畗�U<�)l�����)αO����e�&a/�cI?X�1y���y���:��W����!7b;WE�l�%�a��*϶�6�y���@�3����劶�h 9I>�2������`��~f��G�Y�����zCe��7�閔.�ԃlEt�LtV랅jR�R-lAYP�<�Q�e�+ii��u;��e#���M�Q�
TQ�ʭ:r���@a��𓃰��D�)�Qƶy����rq�tn&��Ul�,B�&���J�k��u%��gw��/�T��+Qz݅��><>��Iw�:�r's4@�E-��@��I��:U>(G)�~���N	'�OH~AZ�����1�f(l]��~�uGQ��ot�Pu�lʈQ�X�e�ؕ�_^�\p9����]�_%����UZ��ޥ�ny�ߌ�sC~n=���$�d�wوZ~�m��C�e�D���QR-�hW����@��'�_��k!N�
�cr����h��A@�	Ƀ��L,[�_�%7�m�*�y�]\w)��RuY��V@�Ҷ,�d��x��Z����"I.޺1�SF��p�I�ҙ�=�mB�l��p�y�f�7Mm���|�^��uN}����ŀ���*���Ӿ�A/����f�AC�t����O����w�����8i�Bbk��oi×L��a���_����_]O�/����:���h���u���_�ht��ԏ&싕'�|+�G9�O�JHyF1P��B�E\uc���<��P^^��� ������ݬ��`YI:pb�6��P8��}h� ��f���ୱ��9E��9��}#�����>��Q�5QM�C:�/ZϸQ��%�rk'��6��� �ga��7��p�:J��H.���G'T�9�&��VT�0�ǩ@.��L��m��gm0��e�@�]��4I���k�R�Mr�/be(��eޖeu4m�&<v��I�؎���������t^�^���#��&}&~�B��}���X%q���
\|�m�xG	�]��2(�K*���9 ���.[������X]M��0��Eo��t|�H�h?��`�	T�?v9v��%�Wt��3������T�Бm5��:G+?��h�͔��J9MR��T�2��oY���Z�Ok߅<� I���C�G0�j=q������g}⬷!B^𣆴�[��[�;n~y.ŕ7v���N|��^_�&ezA��d��� ���a���	z�����k��s�\.�n��}�k��38�������T�SPV�W��F�N݊q�o�!��#�Й ��&�_�H�C=�T&RUO@ ,nϖ�7e���#��)����.�zi��3�՘`t��lp�8>�yy퇧���1�`u�E��~y�u�PVH�57�C�"��\+��K�ȝTo��ɉwk�)���D�ba��k
�q,�!�����ǲ��uyiJ,���8�`�n� ��`�|͞�iAR���Ŝ��)�ޖ�'�Υ�a�����`��-�9(>��������В0ن�a���$�Nؗ�j�L���8qiO���z�3 +n�I[�L��lDC���-����dg2�k�{�Kΐ����g�Ԓ���zrni�ƗTG[���P�4h6�1�c������FrVl��S��!��x� ��O}"��
���?�E��a;T%�"�Rӭ���h��ȮF�s���Ƣ pw=|xa}u5�"�r^��K��=_S[l��թ�i���Y����)S�!�"�*��ʇh�>q�0rbaz!���3�>g�.��0`��q���G%��?�E�Ǣ:`_ډ�[���$����8z���(��p��7a���% c9���^·j��[3��=��HE�͋~�����I��)���+��R�fw�'<�ӆ���<�Qr�����e��1�y������`k�с�����+�X��
��$��'H��q#+_���^l�.Y�z�ǴE�m~���	�m���z'"�92u�<��x��X��@�e�3���ff�T�KC��G���u���tV���3k�t�.N3�-Wx|H�0B�_e�zB�-����JCD(d�=mV���"�jъ�a��M5��5x3'�t1D�ٜ)����CՆ��|�#�%����3�qַ_�ܛ�bO2S?}��S$�G�R�BNֹ���[���Us.E���Q�9枒A�H�(�އ�x{_������O��l�l(CG#Eh�~��R�L��	� i<S���Cً(R�;)��LQ�w����G���oK��K��3���j�B�5�r�5#������'��i���k�K^�ܿ(�o����mf�S��Y����P�0�����*)�m0��ǿ⥣��.�RI�:�`Ċ'���u9�Ġ�>p� �eu�4��%��$8u�G���5���""��'�%$j���p�w��{�dF�,]��B�+�+#��ك�Yq�z�t�ٳ�
����hX��k�M��U��57_�? 2�ȯ���� S�@gC�;�z1o���h/��E0���r�/��	ME��Ӌ�8(J�߭��"��<���s�i_�:����z//�X��Ɖ�X'J�� �un�:�PPf���]�6ȹ·+�!ץ�4��V���k�i_�����.�Q��$L�*�(���ޟ�W�)�y6�A��+��o���UsM �Rfy�y2ϊ���#b�ࢻ�2ReO��]��)���Dҝԍ�cu�͎+�(.��z��|���y�O,�c\��m:���^�,�����A����sW9(����SG���,X�^I��q�c�j\x��U��C��$����
#n�T�|z�I���Y8ӟx{��^+��6��+y�
%�"�_��[/�a$`��p���7�B��`X�y_-�T�f�ց��Q)kkBG��@��tϤ	�n��Ȅ���	�0Z� IJ�d��͍]\��@[|�a���s_3�H�8V~>+q�I�'=��h���{S� �!�t�␹c�O��cɖ��Q�������w.Ō^ҍ��N��2�����,�gq��`��߭V�i38zW�h�\�+A�fܾ�k�Zbocdҙdf`�0�)n�lT�
�G���q��*�ҤP�UߊA}m�OˀK)�қߢ/��̧L�utR��Fō��	q�����:	�&�M�&R�mT��'�/,��,�V�F�T$�9�b�Sqӊy �����H��u����|L�ߊ��gg<��ഽŗ��[��#���M�A���&���ب-[��$��"@K�L��(��mv�4� ��,#�AE�Y�X������Ʉ'��G�(')vև�yy�k�x��C�����������ޥL�Uq�֫�is�C�:�&�0���ݹ�4�:f�4���J�قy�FF>�{�����d�^'�dL�܂R[��˅����S�ꍒ���ԋm��Mߐ�����9(#�JԴr��y'բ�ޤ�	��<�����Y�����W;��ZK�)��1��6������z��'ɜ��.G���z���l&1�2��
/����F�UĻj��6�7���u�E�"c{ܨ��"�������,���<���7g��L�*1]���v�}�b����V��C��	��%���Զƫ������i�l���
"2��Xh��8#�%[vD��������<���Nak�O�Z���ő����k���NG���~��D��p�C3s�i73�.x� p7�|1�Ή�|��q��?��9-��ǰ�����e�>�q��#Td��P����t�'T��*�"٨�� ��p�e�/ �`�g}���P�*�r� (l�AIp�RY��^F�*��7��M�����qM�����*˼��)b�UK<��zft�m�?ZH�a�]��P���9Ҧ�m��Tw:�df�]5c/�G��3���*��|lZ�P��B��3���v+<y�c�5[�j�zQ��jk�dH`�ca�W%�B��΀hnW�B���n�Hĳ�WA�=�?�vZ�8a2u����U"u�(�U��-e����[��.�Tc:<q"��B)W���NNJ��G���]�h�O�L����cR ��|��J�Hw&A ��m�,�|��v,�K��#���\�]8A��!��f�eʹb��u�J�p3;���Ɣ�SU5D�ct�=g{��4 �P��߫*zE������~t��|0�E�far�q� #�>vE�"�R��jv��; �wZSj5�����v����'Sf�݃\ �o�6�H�M4:�G�q��*��N�]}�!XA��v�X�UH����Z��BCհk�U��qfk����,���D2ZB\�,̪�;�VBX�_t��!h�ʟ�H��An֯�w�D֎��I���2I��my��N��:�r�ܣ�klX(�,�N�������X�}�O��V��m~�|j|e*SO�'�4�g�i(R�j��rF~4�*�mj&�A���Y��B��)��1�?=��5��Yk���Ve۽C<�S�*"1��f��Vt�T�Sn*]�ϖ�0�"��eOq�~�Mvx�_ގ�`��
&���q�Z�9H&[\�"TH%ڋ��\��R�Q����S\<��䝹�'h�l�{��v�Hb��R!�@�S���/�y�*v=~��'�S�*:P���d~��C;U}�
i��9̯Tx�lˠA���9�y�.��Pu;�������-%�Db�8���Ǣ]��6����x�k���aE:��@�9H:~Uh?�b:QF��Ft��igT�}?�褧/"��8�a��$[Ġ���g�Î;z�1�j�}�S�{�/P�o
��/�#� � ���l+�f/�g*:�'����l�F+ 1�	2<y�#��~��B�Ar'�"��q�m�A����?�ء�_�������,J�����Ϥ���ʸ( �V�Ʀ�\�#uG���R<8z��x��^zUO�o��"zf�w���Q�c�t��TW�s�k��6�Ղ|��YR��K�t7�^��viˣ��>�D���8�]�U�Ɩ�L��)��|gM�0,��59�w/� ާ�]�޳��<�.&t��CS�B�d��~����t�N�>��=�-�I���ǅĲ5oN�-O�^�R�߬}X�uI{�\��Þ�Z������F�|gK�����m�t�^���H��U�5����HZv*_x�g��k�)��#	����ԧ�jO^�Rr��</(��ϖ]D&ҖA3�&�Y8UO���ĳ՜��AD�X<�`~ŧv�B�1JOo||�'�q�}ҙ*1�B�]�:^�n[����ȣ4���L;m���j�՘w��� u�6gP�0V7M����{@w�sX=:�E����f$�8��C8{�i	���
�� �����(p�ū��ߴ�^`[���x��	�&F�1���&�J�z�k��)~ʰ
����17��@}� ��r�w;��N��K�7��	_H�v4��R�G����O��?��fl)+wVۙa6����5���O��*(5�a�č/wT���&]�,�gva8�����.$����P�h�1�	�F��=L��,��$oX,�>����)�����9{��b��\p!`jM�S�tO!`�Е��s��h��-�h��$J����;M����t^�Mm1L����e�fh�MIp�g��5�T:�y}:P)�M!���:X+ح�mP��{$>���JkM�-���P8�vU}K�m�ކ�b�me�qZɖ�Z�>k~�s[`{X�(���4�3�/��3�4�K-R�2R�n����T�&�bX�B\���/ƍ�YQ���+2"m`�ȩ��&o�l|A�������IxKz�/K�O���S)E@j+��EQ�[C��-����`����˽����tֹ�-57���WLl���z�A�~���.?���J�=�|��&���#��Vh����i;%��a�3����#�IMa������V��Cڦ(���>K����ڂst%iB��'Jw��)Mt�G3+��1���ƒ�QG_4��D�=�5�ь^P���2��.�����,Bk��g_k�Lg���I���Ep��1yb�Cwi��Q��a-�|�<�v3�{����Dt@W�dũ\�dՎ~����a�mM����,��n��Iw���O�e9Q�6�W����f�HCp���~r�:�(�_�q�N�eqkc>4�i�O�]��k)�	a~G�P~+o����ǎ'E3�()a�{.m�l'4��m!�l ?JN.,i �B��Q&�>�s�#��GX�Pg�W:�� �oƸ���;�A\G�x�-\�7*�GPxfq�|F蔋�c^��P�x��O@���$�0{Ł���vK�%Hl�Mɘ �|G(�����/4��E��R���Ń�^Rmܲ4t��p!��ֻ6j��]RܥN�Y� R�e�W<ײjj��rT�"Ӛ�Č�I�/���ǁ�gn=�6�@��'��@W�5�Iú<0*5��y2�t&��g�����8�A�}G����~��S+ ى�rJv��ldf��E�����_P�z|\�ʒ	� �
�e�wN�%�y=���'3��=D�1���7��9���Mե��]��Kl�@N�F�]E[��ǲ��hnZa���^�eO��_����k
�$M�HڐBWK��b���Ϯ&�K
'ӵ	��:7��g�6j>��Y�J⺵�d���l3�EĲ���m��Cq�CPȵ:w���[ ,�r`�E��Q�~zۆ}��87�L����6
�>�q�n������հ�@c��`θC��{-n(�d��.���w�`�k��k܄�h�U6ݓ=<��[ ��{�AVN� ��;���~3�[��g�*ɞ%���Y}�gz���hP���K���1��>���������c�[h�,�2/M��ܠ+��k5t9sZ$��#�;�j�o��>�`�Tdi���sQ���o��j0��c7��x���c�}���@1���|��}]ץܩ�: \w���Ǚ�uBĂW���]11�@��`	%�������:�7�It���	&>>�0΍�Ƌ�ɜ�Far�t�[�E��ѓ
+��U��7�0���mȭ�U�d��"��T�~�Z;���k|��y>�]���8G*^�ð{ʵ�v��l��*���'��q^N_ft��@�1�����>�a~�^Ӻ���%��ړNGO� d������?;�ҷ�벘�� SU.���2�Z�ZCf�I�u�>~�(;�� s�:e.��>��K��qKϨ��D�;m�r��!�;��[�����a ��q��P�V)�5р�����nx�7pȜ���;b�����X�1��Q�p�� ��w�O+�
7'���g���	Ƣz��Y�*�CM#HE�Z�$�E��?|Kx��eJtnݼ%�k��D�bS*[l�����_R>�����⿦t[�G�R��/�EHm�-�=)w�`F���� ��OnX9�NLR��
��$$@����:�$=<�o���c������xd�@)���ʱրyk�K��$rN�o}��=ԦFvr��
P���G�J:���`��(�(��j-���y�B_<�n)��p딣�U��ߺ���,F��鈾,m�:9�Q<�,N��Snߺɐ�Z��4�2҂M�E�����L���^_G..Č�����%U7��`����~i��)w���a�k�.Tln�l t�����q�gے�po�Ġ���`�n��v� �M��EF�*�F:��efp����{�6~���3�&�,�(�N��\�^�}��Ү��ʃ�d���c��n��vYH4J$�p�� �R�����RSe��*l����AI���-C��m�s46uhx�ϲ���~D^�����qu	y 5qYh�Ѓ���s�Rݩ�������߲�2`�]��6�X:��B���(�dDW������k���>��Z�I,�!��ÂtZFV�)�	��豭��fX�WÀ�;Cc<ε����AVR���_�EY�?�����sPm|��?�$C߷����!�A �(xU��	7bn�BWN�)]/.r8�� ��	j=�4�� i��e��J�r��^�f��M"�+�o}ea�
?+�;,������[m��A=�w0���}`���㱾K�K���<~�'ob(�2V�\�z�!���o*��.̟�Z�S��<(�+!)��0�����1���b�-#�7&j]�wۓF��h�d��Y���0�e�Uldhw깧H�_��)�܍p!s��U��s��BE#3<vm�ze���y8��#-��V8/�%�K���b�I[|�U��4�T���iÊ����h��ݸ��h���hp��]�p�8N�������PT��E_I+换�m�^E�b0��$=�n�q�חX+��{SZ�z��/G�h2�q0l�4�����9���>n>v�.|'1�rO���<������-�"%��E7���8�`��#��@��G@�˪Ќ��H�2c�eQ�fU�Z�P�瞘����F���'��'l�.�x<��$�[��g����&a)/ �i������������\��|<V���x�>@� ��L}+��xu�Ćm���C��(8�����}&(��9s�XFD�w�����ճ�c��yh�2����� ������N�v���D���y`3�=�@ߎ��~2U��;���M���t!_k8�ʎ�n����uFq<Y�Z�����!Ұ@al/������������F���N.���/�K��ؒ�@�\*��M��dt6�*�km��ݕ�}��P�b������l��S\�����vuJ]����x8(p�fI����)UUK�uG�TFN$:7�ߺ;��p0E5�[��ڱ�b7�4{hg�K&������2H(.E��L��S(&ٴ"�Ƙ�E��Gǀ-�7Det�-���Q�´ �7/�9����D���Wo�N9*�I��G����L��DB�d�VfW��u�i��ay����5���5�4�v&rPd��Կ��;�TJ�v��U���D�ul�إ�&0�R�j�;�_�^�x���[���=�P<���E�E��\�$y>���?�d�|�OE���������:�C�2�@��\�Z�����Kͮ�S6�+��5ʨTZ�p��a<�-Yq��)��c�y��0�53%�t� Q�)��_��<�(W�	,���MdA_����8��m`�� �Mk�:�l:q̙�	�ݳ��>H�L�������؎X���tt����ɟ��x���d_T;uO���d:.=FR����������u�Z�;\k�U䮳Y����蜱~�']T� :��,��CJǁ����Ӯ�9��*����i��ێ]n6��� ʯ7��
���#Z:��xwq�K�$q0O�{ce�t�$Â�9�C�m4����Q�y�lE��ej��$���[Pm|�'I�R��a?G()�qJ�4UKz?Ԟ��u@�wJDY~zZD����R��(�߸g�������/��K�r����X��
	��� ��e���僧�jzl�}@3�2�=�-�ƹ����Et�$?gGx�H c�G"Ê�kު{D$�h�"�k)�tHW����z��ZL���LBp=m���jDa�A�J��G��D�08 �9�ϐV8ø:<������C'��z���	+������;׃�S)��(~0P���p�wDq�Kc���զj����N�8!@���oY�GG�t�� ����(�8����f��Y*�r�ż�f��f�u%3��{T�7��W:&��"O�e�]��U p�#�~Xu��(}��7�:7�A6EI��? ݇5��Ga�3rƖ*�����T�Y�����Hmm�Gβ�F��VJE��<��B�4��C����`
�SF*����5��?ܳ��h�?��i1v4M+B�X�y���e�4?�s��|.4�g�D���
/W��7ר�&7 :��� O��i s�U����[1>�;�^}��J3��X(̍�Z��K];�[�Yn��u�U��zΕ]U2��S��Ĝ�1˧7&ȖR�үf������-��M�TN�3!!�ov������y,�@��s�0	�R���)����ꮪ�*���/�'�O�����ӱ�aߠ�6�0�"���� Y�,���ظK*��3��x7)�eү?%A)X����8s��`TΔ��E_m�}!��;~�\L9�j��Bm��	���fF2�ťs��7��@%�/�R��n��(A�O�;\�V CZ�����L}�A�&-�yoCB��O�U�Eps2��8?>�[��i`��/ �W�]�>��7RGӇ���4Y��yD��	j���i\�u���`� Ȝ���[ӟ���Rh�&	��?BD[l��{L��2א�p\��D.�y��(�_��@�K��f�c�d�I���HQ-|v!�^ei��j���A�:��9��j��l��V��Xl1�l!�a oS`��X"�/}�4H��"�,�n#e'rmtn�m�$�H�
�j-�b�6tj�_:&_D�����75��n�ႜ#���7el��"/T��kid�M7���w �*��3S,�퐬��t�n��!5��A�l�?޳�>XZ�Rh2�W���;>g�]Ϟ%�AϿ�D]#�㇡�)�CW��·�uz������/w+_l�Ǐ�+$�4f
���L��ձ��ܓ�@Z�՘<4�}�o��eXݎib��F�A�;1:�P��%��C.�z�I(պ?q�]�h�<�j����8Wh��.N�,� �o�Y!L�I�^�@y��a�F�����e�UR�l��i�Vߙv��91C�S��D�G�	��9��L��1Tɭ[�Ja ! i��<���������U�����	0q�`Ű�"������^N�d�)�N(�����Q�8�EW���.^�Ĥ����^"[!*�d
��q�}ϡC��Ӳ̯ ���j־� �X#呋��;ø��Q��ܨ2���,�6'��#ao6tS!< �;G #d��M��}�L�������[]ݴӗg�F���) ϫ�e˝�<V?�S�����-�����O&a�
�UTF�?;�ZN�d�)rF\�N�V��q�|�t�6�'��P��i�5o1D���o�}�\�����og��~ffq9��f�e��+U�PcH�^#�X?}=�� 0^�b���C��l�;��IN�`U�D���sW$j�U���D6y�ږ����X*>d-SA����~�MO�Súꏀ���V:�fc�*q�|t2]� �(we~��i\��0fu�`��/Q�z����Z�iip���oR�g��E؀t���RS��Srw��g�+s�-*��� �v]q�2l��@P�l�&C�+�l�1M�S�zr#k �^�V,��c�ʊ������W�a����D���p��k���22���K�P�R�7��-�:�k܎�";���j������Ya�S��dQ1:נ��"!��;��/B0	���S��	���1�Xy�_I᷏�KV�!sac��� *?���x�ZOø���L~�F�h�N�4X�'^�þ�XzB�s�t(S�nW�EAGw#�AY��M<>���`��!??^.ˍHFWcm�%�����d>M��4�\(�Ɍ�>�ZFǿp6���Y�+Szqb���7M��a+�Z�E��N�͌,ݙ����`�7���f���_��?Q�OE��8�d�H���+N[����Z�!�b�pI��¦�$������]k�#�9�ZB[��K��E��Ey eZ�1btuj�s�8�z�LTV�w-y>j��N�B&C �z�[�����v(�ֿ�4�azo�^�$6X'~���f��WѮ��|��
��R:>��͚{V�� m�����:�pN��57��+Iz�8��tm��F&�"S\5
l�Bi�.\�$Yп�>CaF�xf�a���S�(��ɳ�K����v/M*}��g���s�~����@����ϐ��!`�����Lٴdqg
�%ƃ6��u<�aȃ6�+>*1���<۠&?t�m�zJӬ7Q#��}.��ZJnC,�"]�@�D��b9��(I\��D�cC�"m"d}�dl5�x줅-�z����$F���� (nQ��yv�ɼ����)G���H�vy81�+F�!��HLI�H���~�o��,/�f%��5�<cx����l4׊
9U\���@��oiis���v�Ny��"���iCڗq�I�9���ߥ��1�d��l�dx��k�d��H��d�"kC���.T:�7R�S�wNH�a���U��CJ�Y��
�˄̼����k�B��P�W0"�
I_��.᳤2�>�ʹk�a�W;T�q=rZ6���������ލ���0����"@af?Ǝ�܈Of�/1��T��z�14�z��Lz�؆I{�AF1��ï�ܰ7�N�ٻ�%�;��=�כQ��(w(w��s6�����X6iA,r�v?W��ٗ��	}����;q�P��v��p�JB��֒'tD��tox�z�IX��;5&�I�Gw�c\�}�P��E;�w�`¢�Nc�P��x��q�bS.>�s�����ۆ��U~�m<�ʄ���F�i\�K����q?��L�K�b�n-�=����V�GCt�u5~�]�j�m^���RvB0����c*?M��8���J%Ђ��U|q�[U���m�̷[�M�;m2�Z��#����uX�:��<�SXϿ�Y<d�;���ٛx�K6�`	���� �.�ϛ�tN�@3bǭ������Z\���@DQ	�8��K����Ia�����=L����Jv��R�d�OD�'��&w��Yz"3mE?B,-�Жađ܌x>х��[�vU`aud��觵o���?�������W59bi��AZ�C&��(gsm'�-9�DܡxX�z�$+�f�v(���Ny�ZY�����=���m�Uz�`�%"9���e@
��LB=ǧ ���,��뿉d���Y�\$I�k1n0ƢAݾ���ᥪ�~q��3�*P5L
�J��a�=WX����5���a�9~��2;Q��f�*ke�ጚZF�Gr`f]�^��(�=.ѡW���iJ "�_C0��F��%Z��g�{+,��撄-;�P��>|4�}*Q�B͏O��k�346vŵs�.�`Œs���2�$QY��������Z���9/2��_�|��	/�uj'ih�l��v�3�(��D�ѵ�h{h�Y׃�oH:o\Z��w�4�z�(X��l*�v�>n�D�B���c#r �!�h9^���z�������#���!k<I�/������;���s��.U�A�B���l����8��=�Am���Z��sL�i�##O�9,���:}�\������b�8˵M���h�J�8����^_=��,��у#"�&��(�{O���ya41?D�5�s(^�; o���#Fg?#4!pnۅ����]GM��#eb�6X7�9�r��c�;�{�p��_�U�|�T��@I�? ��AE�C(^CH��%�������Ї����m_˕�K0���cΕ�XF���I�LT*
��7�q�~Z�|�t�9�>a&י���Y�{Ɲ��	�{���Z��s[k�u�����-�7|��#������\�j �qe���_nq����i'�����T)�9�lO��q,�`���:�ď&��6K˕aD�n���vP�Y���1��> /[�Q��W�ncpML�]��?�C˷n}���&1�j�Sgܧ-*)�OݴY�u�܂r�Q�.��)��?�r�K�7(^5��-��4�G�-!_�Fq�h���	�E�v/8(
Jע��V��C��A�@Q0�ko�Qw�p��"[&�~-/g#I�5�������Unm��m�i�@��`��>Y�?�R�uxFQ�,E���K( �8&�~�>f/ʛ��Z��܏D�vΔ�o�N~���C'��\k����bB�=	YaAw��OPQA������ho�� tY�N�?�=�Ma4]��Qo�%�W#��s :�Q���]�@
ih5�^j�4���~_��I�k�����R�1��j��K�%�:`���Y�1���{:���n��E�M����w�de����b�[Йa�^`E��@��ˏСt0�Pv�U�l6�P�s���FQ�ī���l�	��_Ę�.���cC�,��ԁ����Ǫ��]�~�ŔZ��Bn�Q#zą >R&s��T
�X�ֳ��lѺ�8&(�mm��٦g��U�}�qj�z\6�=�4���-I-c*��_��:Wf�@#���Z�u��Ҙ-<��q�}%&������|�.�_�.׵����߂ `61�c��,N�51欔��)ZȬ�(;�ՒV�X')J@<k�Z�PcΟ^�õ�- 8��򧄭�%�v��b�P��x�; �Ñ�J�O;��k0�J쵍�2w1R̀�)��J?ZOu|kyr'�ak𤡮��fմEI(��5�$�_�k����H�E��˕/�6��L">k�y_O7aa` Sͥ�ro��0N�,*\�/Ĭ�����g��|lA`�'��Mr�@����J�Ljؠ�;n�5�줏�m���\��<C&Ƽ�XO�U��vo5�ݺ���Zh"�Yh��e�ͮR�r��k:���?���;�i К*ψ/�h�7�8^z��p�ˮ\���#�G��+qe���s��a!��U�ܾ��Q�:F\��L�x��!F�-iVM0�B�������$DG����h�ط	�g�4�c�[T��8i��rU �d#pC���6�o��K�ʇZT�}4�L��[��֬\�@��;H.��ci��S�86���-�웚���ǑW�*�, �0��L���l��b*6l�6i�ű�V�-�2�-VD�
�(�b`i6$r�'��?��Uc�Ϸ!�|�֤��U{�:g�c�b~��m�R��� ǝ�x���;~lB�ɏz���G�'A[����]�������i���o��(��Ĭ��j�F�A�	֞�E��Mu�_����萇[d�	ϒ�N�j��\��'�j��{��\,|oI4���M8��K�luOo�jn���Q�'��i2��RyQ���w���NeO�	U�0Bǖg,���E7CUx����4�N�Y쌍��@�Z��S��������RST��n�����϶���{�m�F�(�Gk��>�T�����Z�nx�w�)�ef�����F��H���]��4��N��<|���pm��]��g����cj���3��Ӆ�.o8H��p���K���r��o� mz(�
J��g�Bq����s���-,1�?pu��_�ۢ��z�
��3RS��p°��((׃�f�����,$K`�R@ʿ���_�xh��&���`�fyޑ^��l���U�'��Q����0����؃+����ηׯ�{���&��%&�(O7	�ў���e���&	�8��U���-"@s�D���?����G��"�,G���o���'�8�!��!���AO` �"�����~4�}p�d@@�vc��iQ��	����8!	J&��l�#��ؒI�G+��UG35���,a���e
:^��f�SY(7�~^D���>�!�B��}�����aB�	�߄.�4�W��w|kqd���*xP,E�޵5+�%�ol��..�(��$JW8�>5���+4�ue��x���i	�08~}a��N���T�Q����9��EʄȒ�-��� ?���u�	c?��G��o4v�+���\�k.��)^�L~%��eU�,�M-�`o�w�VT�2b��QG�.����L��b���;�zW@���������⁔�����5_Zv)���������@�ru�(��+WbC�U�y��+��蘃k�Q= *��*���(�ݍ�%�)-&���4j2�*��~�+K����2��\���� 
 x�(g�dʧ�aB�O�����k�%�{t�&��ǩ���f���ck:�b������˱�Fа�8a���^��'C/�l�B�iD��̀�Ӌ?�mU��I�@��`9��Z^e�a��0��˄�{։��[��i��th+iQUYk��2:�VY�N�=uAÏc5��Fr������*�r�_�4�"{!����)���Ǝ��)v6�I�_����	���tONX�<d-�+Is�yK��|�3S��6�>vj�˛��X��0S*�}��:���2����f��G�֛gAM�خ��:eh�A�,�4���<3�v>�I�R���]��ᐿ�6�5����_���>�F�闳�0/$dȋ�j��/V�C��|�n���ZR����)dBJ���>y3!�0��OMQ�^��y>�~�#	��j���>���5e��Ksw3�Q��N�s�@�N����oD��UTt3S�6;xۓ+�vy�E�-��n�{�O���OR\w�6;�QY����չ�Е�(hT���c��i{o��7.�8vd-���As*�9�g�`�­�`D��.�|�C�Ӕ�ɥ���W�K��tcx(M;�oP�k%
�n�̋�A�n�~8�����Um�jD�[+^����}���)q���i�1��Jx8�7zPi�a�]O?/�
 t��)���v����Y���f��p��� zd �m�f���W���l�|��߉�_YД��k9Ft�cm��,�7A�0�2�A�=��oj�ϭ6@o�6�l��2��Ƅ� ��	Uⶌ��`�L���T��3�z�ʫ_<�l�궘|7,4��k�䌨�ލ�*L�h��x�FJ�×���?��]w�;�~E�s �5'�;'�s����(��>��[�Bc��R[Ѽ�D��]�$�J�l�-gf��KU;$�r�^����=�$z5�1Tӗ# �kvqN���-�b�lc���&�)����m�5���5������=���b`I1W�M�C�4�7˶M����ŧ���W�˒O:�v�����(D+�#I"P	�B��1do4��-���x\Oo�_0V
_��Z�0���&uT�ѳ:�(��]ft�����H�Y٦<�!�_u��o�gQ1�G�Ur$�q/(���b���3Q��R����Y�r��G�U�#���|C�J��s
��K�-o��E���O��S��kwc$�{��OY��u_�!��A�@���Q�C�"7iX�~���FM��Yy6<|�4�*���s�y��)��#
���Tv	�	h�x�Z����E��
�w�H]黭R�s�ME)&�-lD�V��8
�C�V�
5�g橺�P�q�(hD�!C���aᰭɕ������D�E�	��rp���#��*� �i�d��p�����k�|5����ݠ�D�na���Y��Lɢ�
���m���+|�=鑃��������,sp�v �}>�����V�>�������C����d��%�?љd�u���2)��D��(�jz��ע��c�S�9��x��c�*5�1�SY@�Y�C&y;|o��J��ߝj.U�}�4A��<�&�F����s�O?y"Y �Y��H|��\M%Y^�'GN7�'�dLu�w��q1�z�{��^u�8�o�L�vsq4����B[���V�tḮ2�A}�y���v�6"w�w�#�vٕ����j�e��~4��ರ��ŧ�C��u���{Chr1~6����� �X� X��I��u*4{�p�uP֐_'�I��$}����	��I��'�pM0�u�"�������Y_e|%�0��@��#V�11 Fh�\������,q�!Sޒ4N��0�2���X��m���zB�1������]A�������$����}�y��Qn�T3�-�E�H:�G��e�Ԭ_D:��Z�� ��X�V!2QО��N�xVXX9�Ķ�ҕ��JaD�+�ȟ�$.M�6L�l��%n�2�^��
�L^��hC�{Πe�V��sc�����TV4��;�+F0�P��r�+�Lar�)�:)u_��~ @������Oa"� �+��Y�q��yڡ��\�]�{CA; 
�jqR�`��4ZY9����r�ݵ?�۸}�&N��F��c�6���҇ڮ��K
_@����5R��Ͻz_�_挣���=��ߛ�)����89e��PJ���%#�Q��f�2q�㖒�>6��3�Zz�0(��;�^�k
μ����p�_�V~l�Yэ�&�_٪[��ꔭ� s R�9��cb� H��Y����f%��$�����T,wʗ�����׳�	Ҥ��<��ͧ�VM��L ��6���L}��)n��RP�c�1�K��u��-v�(�R&�����+�4�X͂6��r3�q�7�����(B����a���&f��X���8I$��`�0��@�x�3J�=��;v'Hi3��{�|�\�ޯg !$����4=蚊�C��9i�KjA��ye�<�;��V���8�u�L&r�ذ�FE�M��D�u���Qi/���WO�� ���_�d����蛾U�~��o>+�Πo��'���Q�D\���aCR�W���]����`�mt��J^2�U�N���a�"����^S�ewog�qo#��+������3��h�\�3���X������ݩ.�OhG� pѶ�m�
�QA5��E���;,�=mւ�u$��I>�%-8���e�<m=�=�!?�I�W��x[DcY����hZo��1�~.dr��y�}����nU��eMMi�M@��Z<��G�3O���/%LW��!Ve �쁘���?�%� ӡ�����?�ۥF�	��0O��ݮPp���'��c�ӝ `˻P���nI�*��w	��c�k�Þy��7씳�Ę`��"J+�щf�&c3��œ�cI)g{:�ғ��	 ٗ��-��@�@���6?<�K�r[��R5P��P��j-�:�e~O�3?�ͮ���X;�M��@#t�NR���'�X{�>Sn�]ix����!^��ׂ-�rOr�z#�7s� �EO�Q�j�[�p�=4�8�V�N�M
�Ȭz����@>#�m2�������{�cA��l2S"�blK����f�K]�yg�_�����;�.�]��X:g.�s�{�����>.2�=�SmX��U�t>��.�o�ua�ie�������V!���=��ر�l���Uː\�v���F�2G������U,�X�7����붼�����9�_NhS�9�M/�*�Ql��q�d��0-~%��?j+x�B�*�U�	#�1  5I�5,�o0]ʶ�T����-zz$pׂ�E�֍&^Tan���*�K�T��-+�J¹s��`�`u0�ci�G�1>Ekz��)�Mo9A���2���N�(��<ᲯW�&<�<nK���;1�7T���*��76�@�ӣ`F!!'V�t�$w<�JIf!餁�7S�4���������ܭX��>"���
vyi����mv
���%�z���ZN^�!�����L�#0V�j��S�~w#Zβ.���w��/-W"£��F��_9?\p��<���j�t�'3�m�\�~~��$q���$��DP\�{w�t�*���7�0�HA�xg
q�CV��ӗ����s��Hծ¸B��;�Ғ4"7Ԋ�0����_��r-�)�C>^�ꋞ�TJ%t�E�K&t,�А[���8:m,�i���N��� �A�}]�C93c�Zqs�O`p(��T��Ԋ��O��'��x�5���Q��ǺxUݬ�a����v�����}b����@N����-����-�
�"ǿ�~y�3����`���6�7d����TJ
�����J�\-����IO��z]��Xy~%�?I}	#$q�j�0,ȞX�9�|�t�~lˤJ���U��Q+�E1Jb4���b�(�V�?�Vok���]!ŵ�&��F�u���z�%���牑(R�'!�?D&�j��`�10��-'����P���WD©<��?���B��n��8	R�� [)�a<Op�h��{�N�l@~��|S���f�F�j\��S�E��L߁%waǕ=��ME��Eu*���8��sԑ���A�+TH��il@'��E��	]T�,77<#$��h�b�ь����I�b{���#4� �%H��J�p��C�`h��ƨ��뇖*c�S
i���X�I��9ElSȑh����_|͞����d�Z�x�y�ŵ��	�aTL�qɥ�x̠��S�����'ogeP���`�R��dy�@�]����QC|��������g�����)���t���3J��`�(�L�헠��Ԁ|��M�jُ�,��R��26 G��o�
�]�8t>�s|����:Ǩf�j�X��[+ŏ+GJ��T��ɞjwϗ�3Xu�cuQ��MAu(4��9&-��>*nf�on���2�������i3�/M9ϸɡN�_g�9�!p���jH�K��М�%6Z.i`q�"���s�^ �I���zEmX+H�������͐C���K�ɀ?���d\�LH��B(��|)5���;��6K{�)T.Y�ׁ3�E��/h���9,>&�#�'�{nd�a�ks����Iw�Eqk�`2�S'B[Ō�ȿ��sN�=��f��F�����{s���^�R^�7>����ŗ|F�l!����������!M,�o]P:_Ǭ[y.��h�حL���i�TC:�Z��o��s�a��͙Sh���6�|�fT���Y-2� �?/��CŘ�K�����L=��s�����g�,B,�[�۔UGB�,�q· ���UZ�G&���Oa�S;����W�����΃>���#����NG����Pq7F�n��%X�=,VKO��f_�*m�s84���rD+�)k���C�~F���]���M���z:@��
���q�P� �c�eL��Ɠ��˳X߁�IE�����Kh��z�Ĥ!-BΜ�ɻ*�lY�I�oU�NͨQFS��b�
;�����M5� ,��h��x�XGJ�Q���%�?;s�k`?�2�Y�K���?I��y�F��c��aj�]��������l!���R�\g�{��|����D�M�*/����'��Pd#+�r�<����"'���L`�H�m���*ʎ�uQ�8g���Qr�����6���?:FH�m8�U'���Ř�`o���׍�Lڣ~_A��2��R^�$�M�:_�����׆nK%�82>�e)���+h��-�Q+�T �T�<�/�4��ο#�A'�+��@�\�#�D��Џ���P1��+L�Op�U
�:��g��V�/
�A ,nԞ��I�����P�5�J=n �*��f�L���ʡ&���&�HRN��r=�r�9��&Q��̄�p��4�Oò�D~�P����`��`	
d �s<���ZpQ��U:j�c[�E�����}�x�d�q�@x�r
�)�D$������c�2�~�2"�Eѹ��+���R�A7+���LT�:ʼ��':ޕ>$��fM��謐���lĭ��m�}��e���=2J��t/@���u1ّ��e�Y��u��J�!��V-����&�����r��hq���"�<����3��P!ܕ�ܽ?\J����z%�4y��k�d�b�]:7H�0�E�3��!yu�(��#3dԠȹf��<Ώ�o x��6�Vg*�O��~�\��/�O��.��+q��(?*��qz���P�,�K�F9�͟;��r����f����*h	�{I�U{����]��a�*a��'�X�?��9w��m<v����0v��p�*'�ex�a� ���Zx�����iV��O�ƽi�a]
Q��l�w�G�M�Έy�"��`Bt#Drt�P�����Ƙ��C��j��P����@��"F�JAgXz�*�#I�����{U«L���lUġ5T�z��0�>j�`���0ux��GW�;q�D���8~��J�%5t ��hbP��A2�,M<��N�q("�jtÆu�����w�k�mB�.$]��� ��~�4��bǞ�ѫ،�\���l3A��m0ܸ���y ?鑿j�����.S3Lo�	�JQ��xد��@�+��J�ز�&�t ����H�dewwm���X��c��{L�W���@�i�ik]2�J?h���ҽ����y����������������>g�%h����k�r�sE��Bmٲ�իib��'��@�L�:��jl�q'����!���WѾ����P4)����VL���Y�d��P3�T��w�ᇈ���!�ϒ��~�G�oA�^N_���������S�GL쭍�� o+�<�yd�.�n�'�:"xՓ��8+�h	�L�~� I�nevZM����O*�/r�d��)q�Y!�(a
P}�.�0��E�,����_��nx�*y���y�\m��)�\W�р6ĵB�����?�j�����rײvQ�E.�e��	������/�\�M�0�m��\��2��k�-ޘ�6�3Kl�X���kF�Dcf���w���K��K/j�#5fGB`�Of�F��<_�a\�cN�5jS���C<���'��He�+�v����i�q7ŐT\�:Y�|ʡR}FN�k�#�.4Df�@�v��qZhh����w�4~?��Ria�Dp�l��)�q}A��=P9ݔ!������:.2B������B�閘��c������:H���]xrF�2��� B�8*�GQ���&�V-SAp.�^A���"@��V���7�������'��v\e|�=�M3�ȧ�_�?C�Z���;_��DˡB�3P(�{킅eE�X/�CU\ޮ�
~�<��+a2b.+u�E 
 !�=��^'�h�b�ɯ/��\zp��g5K�4�N��1��V	9Ԭ�ϟn<4D�aq*��28�N���� ���'�:0tT,�b}�'9H�mg��W����pP2ç�X�����b �vc�8��P!�n���v"`+)L�����0Qd���B���j���K���pt?2�R�T��xUE��8���vyL&[�V&�[�UH�&A���>�cc�)�څ�GzO��1	��= ��_ǝw&g�D~������2>\�(��A���%���D�e��wr�V�&�Z�0��|��@��2��}��=f@���
LV�m"X\��4���\Q]~��5�9f��V�4�Wx�o�|��)D`ҿlB�C?� w\�Q��x�V��_�������uPj�*�z�cVo�-v��n�XK"S�#�f<Z�s�wVΝ��HJ��� �F�� �%�!�<H0�)�+S[S��c��Wej�'�@kB�->Mo�k��ӟ�^�\|����Xخ���b�l�E�wru9/�K�H�m�R�}�L�C���9��({�o�E��ku�T��#PH�T���� h!j�}���[@\2��;(N�����#<*|�_j'���X�|~���5	8�+D0����s+|��
�E�����[d�n�|(m�!��*��O�}L~+�h�%��|�|�B��ѓ����ن<��t�<�Z��.�/�~+�R;8�U��#�N>pz�t�&/&؊��@�|51!"G�FT�4_x�3n�VV1�g��
�ɽ3��S�~��ݹ'�:� �L�k�N����y5��N��js.��	u4a���7z��~j�6��jPtr����2���e��(V���g���x�pp'ahE�4�tG�҃��L(�b	I_����r��|����A\Z!\�-�ŕ8�$�q���bc����oU��{�P���D��BO���}����Jc�}�6"3��v��|�L�"�5#Am M��d��W�"<�ټCB4������e��}*�$I�����`��2�(��p��C��]�6F5�I�k�|V/�(��
�Y�Ǵ�aaN�f)Y �>��Xf0�ɞ2�Iu�)1���K������0|/����?M݊Z�##V>����qjé��&{*[�b�q-�
)�	k�dL,�b�>�'Y�N��R˯]�6w�?��ey� ͕���׋I;�z���ٽ������Q���-�@���^{6n�Z���S�q�Ds�y�[t7dR���\l}Ś�6z����at"��=Nt��SC=���x2�Ys-�w��ƴ���ѧ�xZ��P�Y*m�jZ�(�MK\�o��O��y�����ŗ�^� �Ubpաƫ7H7�:kut�5|8�����ܫ�⃔@����÷N�{ zȒ�� >1b�b�,�9	3a���9C��NN�z�c�x_>HHs}%z1D�&�W��a� &R��$��k���--Z��05ib/����$�'󋵣 'xk5Xk),W^d���8�W�ˈ@Ce���<����0ة���b*?A��B���Y[$�i&tc�E�}����z�1"0:t+@{i����[=K�!N��)��+�`�����﹟�ߏ���odٻϾ���`d���*�?�P��$\��6�, �p���߸H��"ȡ��������@�'��`��<0�{oD�aΝ�� �taV�Y�#�^Y�;0�iu���
���@�QEw@N��!ڝ���/<���i�^������p����}n�������o���2��	%�<瑙�*7q4��fu��<�^��,0y���/l���t I���Pੂ�O����Ago���[d�>�ش�D寖�|lE�߇�/v�=R�U��$�(muA�M��	s�%�����c7q{�`���W4Eζ�׮]��m���3�_��ȢD+y�C�!:M@�<�W�˲+OR��=�qx��aP?`z#R��͜��?,�ɌD1���[��6�$�)"��UF�u������M|:�׸���Kb�rD�7w��N�����CZ��YլQ���[ �@+,����W��׻vj䰦f�6�j�RN��F�s�Y�N�l ���P�ι�ۈC��P(���I��?8��|�s�"u{���?�\��j���<��3�����K��8��������g�.��d�u�p��c
e��GC�|�scj��ڡ��%�K�o⻰K�1{S؏}ڎF�2)�U0p]�Kw���]�����%���
ЀëwO�@��a�O*����`s��(�ܯ0����9��]h3LwW�G(�2��.��T�H�_���� ڔq�qC~?I�F6B���1;�����Ebj_	?9�?E$;'E��N�M9۝b�I5v@���ϩ�4�����A\<��>��������p��Uz����d�Bn��ӷ���!U>�wj�Tw����h�wnT2��>pi�>�f��߯�OaV����-�Xd?��`����t2~�w��I���/I�Ά��H�NGM+�߂����2L�˦]婃1���r&��x�xKG�
�/�n�V<X�e�����A�@�����K��+�ۇ�����$��f����;�/�F�5��vȮ�[S�H��k-�#�.>~��.H��@��W�(��y	+��mÃ��!$v=^P�dw�T�@R���=��� v����"�D����g}��J=��"y��`
(�œ���Wtɡ�������39[�y��.�`woJ�I����[uPϙ��Qb�|&	D�u"v��bN�O8Wl�	�:ǣ������y�0*�SX2��K�\A0<��V��@�+%C���nP�4�D���������t�}�7G�P���E��u�֦�KF��V���N�� �z �g�PJ?*(N'�Jp*&8U�+������j���AKG`P��fu��蔈aH���d;s���p��r�)nh��<�����t��"`͟���:L@�2�eq��~�����~��P�l�s��E�T>��^<�˹��Y��kHι�G��u}
�<7)���=$%�J��ƹ��I�ak���1!��������jX���)�1�?^�RxjGz�]�;���k���Mx���J� ���}>���kex��dIXj��h�\��Bc���y�ߦ<�5�3#��j�J1��[���5���<FS̕B����S�g���W��>6�J��z��R|�Ȕ?f��juBPF�B�{`�Z��]�݃��RU|D_o|�cD�w����^ꙍ��G�,E �&��y��%�_σqTUD��.�ӚUoiD�q���:�z��{r�"�]//�q�>ƣ���!�
s���
Bl;~��[8�4�H$�������	���ŗ3t\�@����qZCn]�k���7��6�Se45��Q����l=�ڟ"����'CLgN�ӥ�?�X������Ӡe-|�����r�Oɓ^I��mf��rkW�2���e�bT��Wy*;Y�`��[�Q��=�a��7�B��C����!�]䈄�r��΄5Ú����e�!�B6���Y��wߺ�m��)qi�vT�j:����K��n���/@�W2�����PB��������J٣��+�e���{p#�p�O�?�q��#��8~���TR��ϬI��A*�ou�,<r?�+p���r;bPW�,!��9�[�:��3���N�!I&��osw�%sOr���8�����u�V��4ӗ�˜ˡ��18쉅77�=���W�*dF���ӝ�'��j_WMH<?8E�����qUX��~ן��M�|��Qe"͈*�w�uA����S^1����}4r�!��[�`8��\˟�)j2^S��2�Gk��S���/r�uE(]���7R��dG����~��E<��:<�����_�n���2%8���6s"^��_�`BR��<��U�Y�E^y�_���E�g:Z"�zO��#@o��rC92���{1�P�K��� ��a���h�K�ݲ�IJ���=���Ճ�mOHY�� ��������i�d�C�}��NmW6�	3!�G�"��X�c��� �����
�D�]ȇ,y������4�`\nk�9z#�:��r�<?L�i�ͮr����ҕ�j�	Pq��i:��KF�]������ǜ�n @Ǔ�|�_�1��ܤb�	ng�����֦�g��n�����ʠ����i��e9�X�L�O���\�N�$�%�^/5k���3�FhUhL���>DB�B��!�W���!^�����T%P��Y�:��QΠ���������Q��6�G��A�:wR{��M��e4�L%Jk�{��
`��Ch6J%GѨ*S"gu8a�(����h%0ɾ�q��l�E�[�; ���(Н���q�v����"��&3�3b�T/�����yW��kY���,�=z��TeJ���h�(:�|�s�����j��b��'XXь�1��S��8�H�`$S5��!�j�2t�䜞ɇNC7_�T��<�<�s44^�fb��L	��3N������"�$���+��N�
���s��$ũ����X�OV�,��]HKW~+$�O_4#k(�\Uv"�3;
9���>����K��p��g�X�rhQ�Ÿ#bd�����~i��R��|M��;l��\��^]�u���/IgӁt_�n�f�4.�$켘���Z@��佌���c�~�}F��8��X��?c@�"z�����׬WK�Zmc\���2��k�}Fa��>��z�o}Xb8k�<T�3 }Ct��J4;�d��.M��d�W�PW&FU�2�=�w�A�!^l�^!%>��K�/,�̪�_���1
�gۈ� <ͨ0$�mPDO1��!藊	����W~ɕ�ȑ�u"����BNi�L�3l�qJs �>�A/��-�@�̵s""O�������@�(C��h��2T����G`T��X�����r�ĵ�d�>�ډ����ֆ�o�����.�ѭ6O&}�^TٖTEO� Å\?��{��DUP�R�S(��̓�ep��	ԉUU?�� �z�O
�O~	!8J�kh�#P�����8��H&> �pm��|N��@���QJ������2�s�CL(�14�:�^�$vt��P/�g����|�]m�d��(��t)Bxe��,�C��q%|}�d��ͽ4��2:�5���ĎX����Mȭ�C��[����w/K#b�:+x�c̬���Sϊ�ڮP/��%C�VT� �@|�3�-�k��}��4)�o��Y������ ��I,�b#+�����YT����k�Z�,��;j>t��"Z�8p(6�u�ʩD��Dj2'����I�f�ȴ1b0��c��f�����PI��+@�]���p E�\��n��1�51?�,�/��V��>�xʗ���(̆��I>�gL5a�!�����"�ݩ!����^"9��Hd3�[7t&ԡz����Ybd�=�ԑ������O�>��!Y���I�h)�Y�:�B�Cэs'X��g����u��&����@0�r�{�q����Z�����Z���:�N#�,Hפ'�hP�"�
b���s�ۖ�+_�}�'Q(���}�uO��Ó��Q���Iq��(Y�lͣ�.�l�
�.����K�R��*5��2H��#_�q��>nk �!o掌5!���E�Xm��(3��i8�����Iw�M�э��"�i�i����"}0Z~�U��;ޤ�tFq��P�8��u|���?�Κ��kh]��]�)���,=s٪�	+��rb<�{����!m+ix�K�N���9B�ڌ�t��&�8��2�#���U
�E�&>���(%�Dg���mU�)�-���=�z������%t]������=�ڴ�F�r��0oT����Hw#�:F�a����rČ�,<%��p�<����RO�o{P�aH!�K��0�����x�k>{[�.�9�|�~�7'rNHT��j�}��,I,DJ\�8����u/y�	l�%ҀA;��쭶�.k���^���?���w���ǣq���S���<�/�Z��O�-�d`,Y��jm�C����Ws��	����+����*LnV�`�x���	���r�沁�F�T��"�����i�k2K�تo�נ�ͦ�{@�\ݞO��)�pWl��!�"IM
�-Q��nq�nZ�1��6t�sme�8z�!����v %�a�&��k�eO��Fb��������j��������:�N:�ԛ(��c�����=�<
�S���%���́Cd
�gv��Im�h���7Ze012�U}L�8��\Iҳ{����X~
r�7S? �k�$�a��P'O0pz!��W��V�����l�[z��Z�~Ϙo���VA�z�m��c/�]��^v		��O-�r���OL*������7[�$Q^<{p�T_LŠ�f�>��������7�HY�.,Y�
�0lT!:e��Aޕ�r�����7�usʨ�uP�h���:ט1n�r�E�[,�<(�$
Ŝ�"�<V{p��� ���`%���l�E�T��F(��ѱ3�5��ꮾG���6G1P
1J���܋A��TOu+��%��#\����w�9h��{jԯ�+kā�Q��p�;MH�'և.!l���d���4�Cp>��حzz"t7EƦ}B\�@�O�n�� 2?��s����!�ISE���B�y�E<�ѹ���{�������p���/�����vY����<���@�"~��;��f<B�ZKK��ݖ�G�ӣV8���=�>���=Oi�aS�x 6�eݺ�cO�
���p���O������'XJ�	�?�f�V�ϧjf�e~F܄��Y�4��|�42�Y�t&����M*�S?��';*t��7\����]P�Et|�� ��1"���y�	/F}3 �>rwdd5>���e�qw�s�f����8��*[��`�k���'�ITy̥�3�
�`��UVr�`�M6�w�w��k�֎��xx( ��zs}��?�7'o2����ī�Wu밄���ޘX�=�6�_�����[�'�V� �z$���ҵ$M� ���s(XԊ*��W�uNLd��ş��B=ђYuP�4�"�듟�0>6���v��!-`�)�0�4	"�s�2_�rwB��?��@-u�9ܙ��:W�?�"�mH����L�PGz�ѫ%�� l�e��(Ib�:87��+�B�^6%ˑ"$p�0"�z-Ǯg'��q�)���,������}R�`��w�L��'rf�6�8�,��u�U7��Yϣ�U�[�+�mZ�UP�,��3�V!iTa&�RU�I*p<����������q��h�+�}�1��t�TBd��Z{{QD��S�*(��5�rvC�!8b��/�؊6p)�[H6����� 	���@*��C��J��ə����/���.�΅ ������-�����5y���S��D�-�BQ&T#于�p<	�?N�g�n\��R�4/���Y��i�_��֧���_�`���&�އr���fղL�l�F|�*M���v6G�V�z��(؇��v�l\_B#�)�	�S���S��������/	 �`!���[�U��
�������Y�U�%��Ve��� RAo[����*��}@�+�y_��ۙ|S�FF�F(�pk��\Aǰ9�ޯGC�����-���D�<�N�N0lg�K�10��T��M[jL��Ú������H���ݕ�9�Pz}q��+kB�(~�>s���S|O9�����x�j���TUr�>�+�y�e�h�_���������B4�f�^��	�8G��xR](	2��3��JV��8x�Th]L=۪�9xM��M�4?}���:���va���e���we��
Ǣ�	���uf)d�3p�X�Az���^�j��>����]�]�j+.A�K���v�.��5w�s�!B�OO��|S}�ո�q��9m^]z�g���.��'̩Q�ۯ?�g��n��9t���ag�a|���3�G�� M����/Y0�`͖�a��|���Լ�V�b��D'�(�!����2�P;Uk%�ڂ�u䶢�#�
�?�d�Œ7Q�Q��w����P�RsTɲ#���c����{qAE�
�s�0��'��$ǎ���$V�a�#M���7��>d��;��-CpH=��i;tM��dVu=��I��!��X��F����P.It��ՖNS;G�Yr�6���;�BOڤ��p ����=f�)�:����~z��(�=7��J�	
�� �����J�����_�Uc�x�9�Sf��К��2��4
~h��RmXϵ�[�$9�G�T'^�b� ���eง��f�H:d�u�[�����oҏj�&�'�ޫ�p�\�;l�N	�>�b;���V2H�`�q�kB����3|?�ϻV��#��[+2Z�X���-y1&��G�k����$����_2�a+�:ɶO�Ɨn��Y��w�ěY�����I6�}�/s�{�-B�/������0�Q��c-Μ<<�������7��ݮ�Cʎ�b�"+��@�A_�a�V[�s�x� {��:M�[�/��P�4b��Uu�E�����5Ĕ���R{��cE�����p�W�� w��@כx�\g|v@fI�RZY�
܋�8��k�^���:;{����o�J�dd[c�s!B�AQ/�g)}��	̏�;��;+�y��g[�y*��;r��>��?�����F�q�y�%����]�9�Oϱ"Yl�kǤ[��1�I��q�cv�������\Ӱ2�DE�)�Mu�]��o@y���g�ڱ�������-�/]��v�g�I�#6{/�+@
��q�M��G��"1�d���ŗG*�J��M��PI��;8�Y=J�
ܧ�}�~Hc�����c��T
�nl��])C����IMª�ї2�a-��ox����q��&��S�J���Ԕn�AA]���ឝ�]V�q���?�/�������=������??]�Y��|��x����-�3�ل|����Y����x���\�<���V�%xd�\��?�٭�PqH'ƞ�K�TY[[��E����$'a�}�l�H<YZ��O��ݩ�l^J{�f��@�qH�.� �N:��8#�n��?h��Ȏ�Y���"�͕��?:�2t�)��έ�2i�8��^MW�B�{�#Ȟ���Rԫ�$�|��0g���t�D�X '\�i�ъ����PO�my�S��L�3�p[��P'�ۜ����KN8Xxb�o��Y9�~
nTA�YA!�Gb�i�*`gݵW#��oeG���X������wܻ@�| �3�W�ӗGV�[D�s�SD����ʚ�R��D5���G�^��o�YW��Ԝ��ۉg|��>�>�/�@�Q�:_L��b*-ZzIF���öBV�s%����?V�s4Ewc$`�T�B���0�yL΢>�w���#K��&�_��t <_*	7�ⴓ�K���� �,Ġ E�S��-w~�$�����4�A�����iT����f��0�>��i�]�4�<llK�͎�O�g��k�3�ޙY�ѧ� 5Źo�l�/a��
������p�4�x��T�)�k����/8�[���,ch{~�f~�� ��|x��0J��{�WI�7�.Cվ�t�^�wg�V�Q\�ܼ�O���#�e��F���:b��O�n��ʟ��5�#L�����)�U���7���⋐H�>=zjղ����,� ˒�j_���c�H>
B���D�ۊ3?���E�0�ËH�̋�%�і�	�-1�,�q��+�*;��~����π���sO��74��9�:�2j�KP.˻���7w�}
@�,M�8�-|!ڍQ�>.N�.ߛI��-$Z��&��X�Sh�Bth��^k0G.h�|�M�2��h���Cg�k.-R�~;�z���JI�6I�C �6A��^I�h�ȅ�y�\'�+�$2�dD�f�~�L�������l��%o�'�w/nS/�Qb�f���B�@ξ[hpf�=0¥?�Yv�%��-x �]��}��K03�r�yr��m�e-���ѫ���rdM^Zt'�+4�jAʯ��	�68Fش�:d�!�Nb4��S٫;��J�6n2o�X�@��<_m�p��m�^.��[ߤ�&GL5T��)\B�)4v�\�q.[������č��J��CVj\����|v��֬������DN���=���W�BI��O�J��S,����Jg��TD���Z#�h��V���L�]�V]C��b�튂��`{g�\[��E�#� �n�\��r�T1/s�
�C�D�\!
&����E#�I��D��+�|RUK
hI��>,fn�WK�\�G���bϒù�r(�N^�7���wI��B�J��ӷ��X���G��>�C�_��H�[��^C$H�˩�z��Q�I*H /B���/��6�������]�&�q�i0'Si�7I�n<�v�����&��,�Y~*��HO�I.�1L����Ъ���ﾰ��B��y�}W�{ �j�;$j��}`֙�86u��uR.��FD��X�v�3�.�0����ʻ6���/'W��>�g�it���K��hT/��Y�N�4l�Ӫ�3jg�9��̛^�9D�{�Ӫ��$��a�"�ۣR@#��~������� w�[�[��*��'�3���Y;S�y �)��liC�y��� �cv��X��ey�:%�0J���=!�8
R��r�������c��g���cy2L���� �<2MZّ�&�Ó�6�ݠ��������I�c�.[a��!�U͙�� �3s�D�F~��;��oa�]��z2Q-����$��*�s]���vNƭ��ij=���f@^���L��7`�y�E��P�9FxN�+�і�Sa�	�F�v�!�G?�]Ȅ��zΈ�O�w��KFG�̎�WS���P�X�\�c�������9P���l�L'ʊ޿.Q���"��=�y�!5\�XOK��m����v)7d�F��?�Nu����Q� .���C�^2�3�����rs�)��ԡ�[	_p����*��J�|�'�H�B{.���Jo.cN�`�&)��3������Uj�6�p�`L��`݋c;0ڋb�m�%h;6a���׀��s$t�Q��-%�T�mW���ԵMR[�SD�!���r�L��Ȉ��������Cvw� hV����B.��rXC<��������$�S��<�����(S~>.��,�IǗ�Q�۽]��@̣���/�e�x�:�G� ���������늎�m�)ܱ��J,��+E���5�l��H����דΥ���.���N�f0�C(�VUO��-���V�(����/�2�O�}�ζ�������_�rᚲ��nk�.J�J�	�SW'0˖S�~�wi����+}�����3�4��c�|'�*��Df�ND_�8,Hޢ�~�TT��ND20� Ǌ��<�����Q�6��2��r�-�>�?�Û�i0N#�WG�B.x��+~똯�Ahe����z���N�C����b��*�Ğ�b�^�� `2�C6G wR��~Ư�����bw31`�Q�ܫ 	*�=���T#�Z?��U�"�[a���d��ӦI$�a���A[g���<\c�X�������$wD5헖%HAzl�7Ȝ���u\C?�l:�����W�g�~�#g�u�����Et��*Xr�}������GD�R��q�C7����r}w	�Y���]_?�
a}��묰'�c%�SY�;z~_�3mꈽ���AK1�IXrQ. �jht��!�E���ky$�]��Qy�9�{�&��UG฻9�hf.��]�]�� �}%%㶖��_!���;Z箹�+%��~nn�L�>�F���(),��++ �y��-�îG������p���_�oښR�^�g�g:�'����1x�f�F�4��ei&H֊�a[����A��F\��u,|�j�����J�\��J�;��j�OVD�.y���g�n%
Ĳ.1/L�o��O�j[\s��kx�H�[]@���ݱ��f�����U/�=��;G�c�]����] #�ܐ_�	)�������4/�1e|���G�ov;�s+|7��,jX}�m�;0}�O��ݘЕ(�?�ɖ�sO�*�̆5k^�鮴x�=g�K��E�3�_'�v�$Ư��b�S�1"[u%9S(��Ao��螕�׫��d�s�E 60�AK��1��3��޺봎���������畵"@��Č@����bC�Oh
iуm:��B��mݟ��Mݑ�f�Y�mژ�C�^-%Pr!�v5Gp��3��x��	 �߮� (�\�֘����Kݨ�ҙ���p�l>��d��C �������� f��DL�!����˰)X��~�jzv�)�:�9f����5`3�q&��@�@%���qW{c�a�#��[��*��c�F�U�vm~AP����z����\�8�`��:>U����U1�t�w�C.t�������Vԟ`)�r�qn�/�NCH�4|�2�PKr'Ή������G���6,Q\��,(��.�'h� V�e���I>;��>��<](�=�>ɡ�+v22��5��]3>�����X&�w�c R�9�J�rM#`��5H��w�1�?��a��A:�h�neV��N�_�Q5��Ks�3)��J5==�V�"	�!����SI=�c6]�9�;o���e��u�)�Gg��\CW�����������f�pLÖ�]r���O=y�R�^�oɁ:j�զ�c��fK|�˒Fnޡ���>{Y�byB�ʒ��^C�'_qo!q��-��M���|�H��L�34��0�ǲ��!�����OhZB4��t�+�	_e�SՔ+dV@xt<��i]� ��vi���!�f�n�q_p��������?p�~�>kH��
k��{����x��^f<ax�����m*
��Hӂ�^0��y�����d�c�Ep ����?�n�r��tg����N W�[�Z���=p���/E��
�w���jG������e6mW����G����|u�]�y�I�*��/�|Z�L�V�N��ٿ�zQӇ�<�uCߚ'�NZ���t�T���W�:��=`o��[r%��Ό��'�ѧj����o���;�ɱŐ�K�/�*Q}�g�d�����f�J�� dN.v�a�֛׊%���:]��M?���ZIZ���C��#Ұ�t�{& k��ϥm��:F�n<.�n ���%Cԫ1���X��ߚ�e�j�$�������ke��^����FD:�/��� ��xʏ��Iꗖ����I�������Qn�yB� ���P���
=�>\�A�4y���K/���Tc����b5*��.C��t�X7�=\`)B=������\v`�o���jP��"�ի���em�f�A>���o��W�]*�G ��	$����јC>u�_�E< ��G���΀��\���s<�
��bi�Ly�� �L�.�?q�x��QS",b��r���,D2�9����2��Y�6��	�4K��_�4��W��dA��3����:x�]�p��d���o�W�g�LSy��>|�J�V,f兊����*I�E�q�t]yO���z)��=C�iJ1��J�A��Z����{���7V�_��i"�%r�|�H�l=1���TQa�]�0\�hl3���RQ�hG�+�5�=j�kԜ���v>8HvH�9�pn�{()�̅GS�~�全���	�C���O���?pB�@��p̰�J���(h�AH(�"�I|�5�Ǉ��o`��ҭ��pi�/�^��g2���QL�o>���-�&#����L?����V�{�c�j�x���9mU������ ��xL�%i�
� �ϊB��G��`�q�ȫ���
���)���(������8�_���\#���]e6�-7�v�K�89[�"g޿�|׆Z?�įƼ��)bs޿��@q��d���D`C�1�21%�RA#Y���;!��u�r�BfGfNH�e��H��(x��X�ٗU�) �(��[�LE�z�U��-��b��
�W�kٻ4����1
J�(u8�gB;�
Yy�i�����~2��v��&]^��lY6��Mc���5�\���\��[�/f�:������� z�	����ܕ��M�gJE�����i(���{l��k��;�71��]�4n�J?�S]�����tn��3��P��z3$�{7O���u��b�}��gCO�.��Z�5���	����t	��CwȀtc�)�d����'���Ɓ��f���vA ��� �I������y4e��˽�Z�Z� �����AO�6ŷ׈��|�
2B� �cy�;�-Y�z��6�=X�Bq�΅]��k��Bӫ�wpu�70
����v�䰵���sL��[=?��w�96ۿ�Q���\��nc�Z����EGz���qE5�miIP^�� g�L*�����ʗ�B	brC����	�i3������e�
An��o����t�cz�%)��{����5\�Z}��oC����W�%U�&,��N��!3���C� 8��x$��|��hnx���t
;ײ�$*D��K	ơ�l	`��R_ �&d�_[O���?B��������kP�f��G7ܝAL���X�z�U���ފ��e
L�f�0�=*Ӷ��rp3�1������/UO��j�]	��2�4)p�pA��w�<2~�m���,��F�jL�+���k�f̷k`�0�ˊ&}9����?���i�g�RR��^��a�����O�{�SGo�`�7���� ο�N��
��������u餙� �ݝK�,�h�ֲ[�"�'i���5.k�<&�^�X(���k�8���h�4�����4���׎o�CN�*�p�_�'��!� �l1_���n��οtpD(�� ��I�b��tO���ZK��n^�]�>Qk�8 ���E��$x!��Q�V�8D��NJ��)#�}6߳�w|�Ka��o�$b�*��3q�	��e��,MŋpcvB��|H�r�UĽ?��A�������o�2ϒ�p��{34A���+���~!&��~�Z�U?K����#@d�`C; ��s[r���n
�n+s�q�����KkH[�뉙*��/�d)&zL͒~b1�����#�Q2w-<��]a���:w�V���WΙ<y�Fs�(�`ĭ�= ��>4��˓U�5 ���Q ����W�N3�g���n�{��Zg�;��ѣe���&lP��G���p��{O'���Sma�<�1z:?�c��|�tly�i*9�+�Đk.�P��SK�O�D�z�ToS�\9��@�z\��ʙ��	'M���R�+=}n���cZt��p���@��=B��(3��Y��\�
�L�`.���D�!�&m`���c�QB����N�k����H�f� )����	�՟h����
:���(��2�b�L�􅶡������,f�n:F�y��8��1�̐�)�}�$ԩڠ�#I���5a+����Nڟ!\�Zڐ�i��#RKE��#��x��~NE���zG..;���f���L3�%DTq�B�	Dc��&�"a���C�<HT����"zC�R�B��Ig+�\�	�!����.� �����A�beݨ__�Qk����Z��e������	�:q��n%5�a�9^�Z�e�'�B;�3A�n�d�J��c��h�����%m��*�C������X��@y��8X�yX^�|.V`��h�45א�EdE �o�iH���#P�?o�<M�V�i�KY6��x�b��Z&�%�t!#Uѐqۜ��L��]f��4ֿ�%�1�'M��*��k�<��Ϩ6O%l�ݨ׫&�%��?�/�`��������k��s��q{B{u�D\(�m�K���)�w�#�U����Q��u�ٗ�ܫ\s�&��T*;�[�xc�>�x�֝
�vI�G��M��֭�3��e��دڎ�Dy嶃M�k,E��,i+�;i�'Pd8�M���È��fc�����|�웓���`���_+s^��}O����ԇ?�H���1�AI��4���p����I�8-�8�(���s���&+�=�)�Ik����cNM<��AA����\�r���$��Gy���3�p��§n��{jB#���
���UŹ���e�BV	# ����+7)�2�÷�VaX} Ͼ�]�%k)`�+��G��Z9��۷�u��\��1zt�������V��lU�<l<	{7i�<>r|�7�ts�Hc����U'��������
�������n��>$]�C�������?.�%$]�?^�� �?k��wO��F�u��R�u����JEnǧh��������͚E�s��0��\s���ԉf�7������"9����3l��{Jn2�Î]J6s"-��4�BZ�c tXCl��[���x��8�ڡ�;5����7K��t	���@��k�:Abώ&|�O�s�B�<�C(3��z�4���I��K�F3��h ������\
cSHi�Ì���3�)Ew0�v�n9c�����6�6"�s���>��3�F��q�?�W
&�\s[:�O�	e����y�X{�X>��4M��Fj�ɥ�(n�N|�������v��Z0��l��H����N�>S�e��x����M�;��PR~W��_SbY���~9�'��6�#���
�I�eQeB�76pF��]0��
�U�=Xg�����I����.�R��qvS�-9B���iЧd�4	Z�Z�͸q�����_�b��T��\�6�nok���po���G�#��N����H@0���	�:����?�袧�X3(���r�ə�T5�_� zQ�ئ���l�5�`����C��:�#]ݷ�~d�Jj�-����݌plGz< I��V:

t�|�GH!P1�֘�Q��b*]�zH�Ԯ��1Nk������
 �;+�VEw�����O�7�0a�[��V���<���+��D���S���[N��N�^�υ\bbk"?T.�]��(�C'5���R�	���"���i�jqP�YU 
�؇Ǥ���d�c�~�DG~�4?��??vq�H�f���N>��C0h�M#��1�U��	��v���<�Op�"�(m���XB�OV�CRn�T�W������;��?a��J���$?�M��:�R�V�=(��>bj^>in=IP�� �=v\���6��%a�l�[n����1El�V[V˄�OaŚ��ٛ|q�g��1Y��ژ����-ma��R��*���Z�~h� �5���J��=��h������h���,]-���1aj�cǼ!o�_ԥ��c� ���P�	�C0�8�[�t��I����&R�z�2�v���>�ů���d7J��A{��!��)�\o�3A��+�=�(Z��[m�ㇺ8ʽ<vM�	���"{�Sj�����]�%��$!�m�OWC�z�q���>�� �w�<p'v0BW�]I�ҸHh[�V$��Cb��f�ed��_$ l����"�Y���O�r������,k�6����t����P��{������nYXLw��G�g�m����a���	����A7>����c�a�H��o��������l�[�l�?� �o�5�����/�?��ֽͲ) ���P~�WŬG��;_+��Btx[BvLѡ2K������`�Ŧ#k��L6��g��>��i���c��T5_���^/�/��,�EL7a8�OX��J�;
�Mcl��TNb�V��9L�Zh5\�l+��c�[�O �n|�R�b��/�֘�=�0��(�5t[(���|�/���8�n*G3��f)�h�bjկ� ��E_� U/���۽�8
���Q�~��E�)�S���ؒk�� �)�>�;R8����ɀ�0�����X��ʅ��������a��I�h����'�ZA=��y�X$�Y�!&�H��\����^8�X����#��ٯv�s�I�����CP��&����$��!�K"|;iop秂I�2ӟM���-p�����-�ߎJv���?�����\�>�T�/^�7��$�9Sbv��ɡv�����Q�?���"��	6z�l�c���b»= Z۵�/��/�{p� ��\�L"�JEae�4J�7�3�&��,�})�Q�ʬ�8{X*bۥs(M>�"���5�bs��F9i�yyJ�Ɓ���2�k���[�g�+4��(@8Ą���=?�Q���3;�2�J[u�y�JIaք�W �u���@x��9.�|��f���t,�FYmdZ?œ7'I�ŵ�-m�Z����2z6y�� l���[WtQ��塥B}8�Ol-���W9��eOp���b1���P�({��}�{C(۽;I����Y���/v�	�sO�QeU>�Y�NJ��1�frгB�A�q��ؑ[��7$?�2��7#�#Qr��F��GW��!�:v���H��i!�D�m�kE��O�!��_G�`��iu�Be�ewM�+�%�^�c�D��MEM!����"�#�G�Y��F���)��w�l_DV��G�7E˰y�|Ar�/Z8�������%���\R�B��()�w�b���"�d��m-�����������_;�τe]~?��H+�*c�ѷ�%F��GYo&�ߓ  �3 �0`����P	�����%�:�?��x�BZb���X���"��;o_����2a7�42��p������0 �c�љ8�j/�k�ƥ;�pY"�D/K$h�@����~p��{j�U��Ĳ=�%��$�S4����OQL�3�xuB�k��0Pusv�/z6A�E��yڧ]��w�/�����W��V���>�܏S������,�؇��)��.��mI��S^*��ʍ�x�S�Q�������ZR���k�F����`�{�:�Шk,hМ¦jR=;x���,91]�5�u$��f���w�����et��ԟ�g���mF6���i�Rܸ,ݖ� ���"�Kk�O�Q��t�zo&�՝y#����pE�❧�-=%*]` �������lC�ܴ���_l��i
g��[ l��b�]�>]�쯨����ZJ��y�w)OQ�s���z�-��������g�w�_�������M�������*:�7�W��Dh�>������W�]]��Xn�Vm=Cټt>7�ĢD8��o�`N@��T�n���TuH����KC�����YQ�a�:��ɰ��謁xLُ!��s��/ �b�7�� n��j���ɻ?�1���抌(���gR�b�^ԛ��1�pK^�]b��̈́jv/����(~8��R_e�lL���A����Ӻ����-{�T���Jh\�"��@6F��c����}�L��L�ŐF��l9("���������ʴ7�=9�I�������M�F��?�O�z�c��S0d�쐑�c��T�3�`�ҷ�9��k*Ge�B�*�sA#؅#*75����������ã���Pހ
/���ڵy�W=�}����I�"<�?���h��c�s�����*�֊uh�T��s�_��C	� \|�uM�,�%�0\7��fH��n��{e�H��I�h��c� =�{T���<�f����M����
���9+��[$��K7Kd�dz�OHh�~M#K�&��<:� ��n NJVZu�y�f��UC�t$�V,8M�~X>k}
��,��La���bN!
8 A��۾�1�ذgJ���\4iU�\��Ou!���1�%R<��dG��V�:�4
6�_��A�Դx��Ǔ���Ybr:���k��t�r�N��j5��"RX�L.���k��_H�	��S�x8F��$cx�D����8t_�L�(d�)Z�"�W�wgw��Gw|�QC�ő�C���Mj��C�DL�i��X��
M~e�9
6q��q"��A��2�K=���7YW5ᧁʷ��^�"UsG���M�rHL2�i���gL��3�R
q�Bә�0�dW������)�8��*�z�B����/�iq�*�˸�l �ޕlA��w`�w�&��Ԟ��8�τL����M_4�=�/���>���a�_�vy���(��S�������%�#C���h�X�l�+�|�>��W��/�#�u����:�| �e^��;��� � ��U5/��[��=�C'D�aԢ1�����ܪ_�Y�������k+��@��PJ������B�D�Fd�,�<��5�BK��ksFZ�<�0W-ʴ��;G^�b
g��Y�0����n{�ceӹ �r��@6uL����ĺb���'�%�B>��Rs)��H���r�E^8@[�c�>涩t�[�8�2�l���0�-��|�Y���+pw$��v;:Ĳ�9�����`͝KV���M���Y
r42����~�j�v_����_(��5���.�b�h�P���Z`̷̹eqe��aJZ�y�`�!@a�;�e޻o���1�Jb �O�EgM�"����dl��H1��8�ѭH��X���j[�����6�F�K��9���	,�>��(~�\R�У6���B���V��+2�35z��n��^\���z
:�'�a�N����T	�L	�)�
��ޜ��퉥G0!�/�N�8�^"h�+�����L�R^fp�u���5W=����:x�����К1�q��;�U����2N���p<��{r�`7h����������稐;&�	L�9#��#����!��\-����>:���)����e�m�]*�=*3hP�z2yq~�Զ�G1؇���������E@�xy��zƆ�1h�H��(,W�#�9w
FW1.��z{����~?͂�
Ys�-W�9jy�
�R������e?ؿ�kY��[��{	�:;H�#}�'0��h����Q)�1���:���mv�t���K�tg]^D�L�7+BI��N�FɩZ2�8&��#��ԋ��['/��1p-��"����6t﷜_?����Z�_�����]�Sg���+���%��6e׬��MAN��F����,����'d�a��}�SV�be��hQ�(��u���y|�r*���gd���FS�z}=O�H�0y �h�i�bc�\�g)�~�Z��A������F������'��L�ީ��l�^�J�d}��b�W?;����4kv��B�}Oi	��>Kǂk[��8Z+���[S2Nm ��b�%�(��xK���j�2�gk�Jq�	j\���1uNFW�C�@��E�:��Y�ߛT5��)�T�6#e+���f�L*S��.�-b������s��$������b�lJ���g��h�%z��R\Y>(�BnW0���N�hw�b%p1!��t��u��>_�w��T��.ց�H1~�G�M%�$����ԇn���^^tφ��i��H�]6�?�Ҥ?���G���h�Ǳf6�6~�r�P߽����q&�FJZ��[s���yq��e.H�����Ĵ�d_�+�I���21\
Moji��R��է�c��a��jzm�R��a��4l=?W�e���P5�K���5VNqأն�ے��Z�� �S�/Q�BM1�h�m�!~��:*}��!A�0�ՍM+�F&�j�2�v��\z�Z�n�u?��cE�,P9L�M�N��h���c�-��.Z�T8!�BmT��=mܷ�mm�@o�KM�0�FX��9^Ns��w���]_>���1F��w���˙y��Ǿ�ӫ�#�s��?�9kJ�DP��utOOM��ӫg�
�4��H��֫z.�� ƃ�"���;@m�q����\(�WPW6��K���'̯�+��>�`_��i�S�dlp�$<7Z٠��Ri��*.�ɭ�ߖH=>3�ݛR����F�*�G�&�YNpO��9�x������[	�S][|{�JK]ޔ��A%�`B8k(R���tt���[�43?_>v���<{����ĳ<�Tm��%����
�9\�~�.�ee<Oo`Ex��v@�FK���!#5��J�E���7��8(�/�G7}��w��q�he��q%c��t��5���;K����F�Y���@V&Thf���u��4��exK'�/�ʬ>��..�c ME�S�2�{e�zy�,	i@�6�l�h2N��l"g�gV Z�܆���;{���4^�8�X�\|�y��ٲG�W����.�}6,�ߦ?�]�8t*�-���x�EַX��O�J�ۢo�9	yY�R�rG*f��
r$�E9���U���uB�c��G' �C�G�L�W�^k�������fN�bf�QR%��8/u�ܜ�j�OhA����z�-W���9��v���1�!nnR��O���c5E�2�"�������ǔ�
U�#�MP���I�ٔŴ��3�BG��)��t9o��������G����+�h2�&�t���A�\�瀊���̣3B����@�J%)b�L�[�=�3���'�6Mjf�"�?q�;%�<{��3�ޙ�qTώ׋�8K��C��#�J?#jM����A�!�|��$���@�\f����kI���a��F�b��_���=O BH+i%_��1wm��
J�ע�푹r�zs��!��`���`7�����M�2~ق`���Ww�B_,��60K�S[=R��0�k�V�`4�o��zN�]�4��*��&���Ѻk�R���:��8��&�sP�@c���_�h\�
����rNF���p��ϙ-ӺB���x�=��
��⚤�&,5��7.���7���l��3��ݓjgL��r��aE1�:����N�2h��$:�pfå&U衋���)���=*͘�B��߂h�yE��<��V�za� ����I�nӘ0b�Z���SR���o�$��g�)��kN�fa|��<��R,�Ւl��e�6��\�F��=c��2?a���|K�^~b��n�N*����-Oh��݂����Ic�V'Q$V\sQ����_;���J��d�w�5`+�&�j��ȁ��~>f��������=?k���kq�Lq�bFh��n0DF�����v96�ǿ��ʘh����E5Q�Y"k��I�|����:qN|���~��b�}.!��R)�xQzp6\J"(��RITH�'�[ϳZ����H^ ���~t)\��(ؘz6ue�,������K�W>���[EA��J����H(��]:���?�'M̹��)32�JTx�qN��R�W%4��9�ZI���BcS���ΉW�ۢ}٫��d�~����<K��ج����\�pH��7�����څ�e�d(�Dy3<m��wOu`�9�ʸ����7B$/����$᱊��UG�s�����',�m�����q��k��C�#�J.�L]�-��4$ގ�j$�S�g7tV�8�Z�$�-��z�ɥ�u�*0pBeC��?}|�a����h����p�9�;�&��L<��^������e����h	�|;;��ӎ���|%/:�-3��x"~�"��&1�R�ڔ�#n�W �z����3\���EX�n�=�*�&V��r�Cj���ri��	��[��綠 [�Co?��%��!QB2c��?6����>��W ��k/L����[�K�(2#���f�J�]Z�>���[Y�͘䑛�(���_��թ޽���(��n���Y���w\ÈZ��-$H�L3�������~����i�v^�&�%�!������Q}�Ў��s5­�cw�~�wa1�HW�Nv4oM@j�jn;m�Wp}�����2��Q��#�k��`i�l�_%�D^��*���I�%�U2�wH�R���l8FO�0���_�� �?FԮ7c��#4dl�C�\�w�f��* T&(w�58!t��݌S�Q`�O�äO#7����jCv���:��'X_�$��=�v<$�%��7i�Q�8�s�}��2[���_��"p��<���(������%�F��l�ע�&��	!���rF�E�)�8�WKL�}�}�&^�D���%T�3��{�
�D1�,���֙��#]euJ�>�To��k͍q�/&�6e���=���8�QRc,�>�`D~��ע�h{ߞ��3�!� �w�y1QkN�U�/������N[���;_ʵ�;�@�Do㸅i�BSed����yg�A�~cL5������Uf[��9��>P���g)8��%��A�q�|��G'��a�<����$� z�N=r�f���K���;Oai�pXI�TKJ��gve]��-�#h ʉ�$�{�j�ᢩ �O�Fۂf��y��~��?��C*������]�Z���z�6d���ָ6��z����%΋pDP��)lo:�Vp�㝚+Q��>�9�Y�nP�8���o�7گ�U��9c��;��7�8j\�s�1n��w.c3Bo{,��+����y��I��)*W6:K�$,� 
D|Nc���E�t09����p ��%YeG5)�~	�4Fa���su���ö�ũ�o�c��K�'��NT�>G}J�n�d�'�`�Gḋ�:�m���{�K<_��(S0:�\���P.�ǎ�?�4p�,���pe��Ge��jLG}Z8�0b��*ZD>����P,X*ޔ�c��Z��@��=k	,�%(�(�rٔ��a`���_[T7�tk����k,�C�������ϧ��2��s>v�B��0.G�H�J�z�K��`�={��#ɞ,?x�)"�2#pI�m} �!��cO��X��\��6�=��(TQgMh���(F�w�����֐��R��ɦh� c�l&�tw�u-�fXIxq+��B�@�K:�B6�?�����	+d5R���z#P�-��N�S��������x�w��M���G2V<N���{�o6w3
(�?���;P�o�m������(¸��$�e���ʦ�����4�K;̅�"k�7 ѓ�,�e��v�5b^zs(ϥ��mQ.��C��� ��Ġ�r�{I�Ba�M�:��@K�C�'�L���fP��n�kO*K�8�mo�V7��	�b���zy?e��B�r|4Ŧ	��SBXC�z�e��p|������]~_ĺr��g�g���8M���Ir�<d㰆'Տ�zu:E)ej�F+7ϸ Bt�C�Sd��b��ZIVC1��
�X5�q%MZ�k訧�S��4�m ]�̹��	�}I����-�1���#H��غ�a��jᵇkw*�j�=-D���l��*p�"�w��\}����֗m�\��.��K�]�9J�P �Ks��.*Y7��a����b{�P�d�S��v`�@�zuU��DrP�����g��$�8�@���w�օN<h�"3�ԣ�T)O;gz�/ue� ���U���N����.M��-�`hsOW_jWc�5 _�����a&5)D훗y!&���([�q{�<c??�Ƽ��3l�
� �PJ�k�h�O�b�c��Z��,6�`�
��dn�gUh�?�s����6�'pD��K_�n[�fl�c�1�FzMu�w�+��uLV����䕛U4r���s�4��W
�G�;����(�����J?��҄P�׮����՚�[5M|��'�)h��9�xۘ��;��D f��,��u�.���p0�VSRēMPbU�����*6����vhR_8A��zi�^S������ �<Lc`��7�.$5>4�rm�ן���Y7�(�:I��j�\��΍��1
�(�xd.����-H��z� ��P���E=y�9�o�j�O!ǧ��e-���Su~@6���(������*�zcL�;�F�p �?+��Xm�
�9�=�Fܽf}E�{88g��md^���	�a(̅˾����pJ�Y	�s�5��_�l$~/��~�a}N[�3�$��ף��.��(���[�XL`'��9��8�P����D%t�Xa��>6��M��ɽ���s�^m5'h]�i�V��+�"��3�fP���][��ꪫ�� ����9�<���zF:K�ڍ��@	��#�i1�X�')lH5s� ����HrA�������	z��C©,p]��#{��ݎ��^��!�86���+U���,�ن���D;��R�w7��n͢X��B�Rg�d<�@�8lj��#Ec���� _l ĦV��,�h@�w���+z�Σq`Lp��FMf@�voϙ�k}�׏�}��o�
��~��½����u01+V,a���� �u` �Ĭa,>�r�G�G� ��6�_���)of��ޓCu�j���-�_�x�U�j:�~F���\\I�,�ߺȳ(�}���ъ]���-ÒrW:p��� �r������J�̰Z��݊�s��|���� �(O@��Ϛ$���j�7�4�D���Gf�K���1YA\�[bó��2"ЕUr��S�;A�iV��Jw���$��U�7�ߥ*���B��Fc>1�#�D�����U-1|�� ������+߆g^��h�F[̃�{����Ŧ;�����=��̈�(���ciٸ{��o�#m��$��3_Ή2E�d'���l�K ����/���y��+��q✵^L�����?�eR&��QW/̹�;�-�g'��z}��L+KÄfI�
1��*��54�3/5x_��������Z���kZ�<Bg�s����r�އK	�Ia���SnbL��́�ʠ|�w_�E��M���.�^	G]pWle ��Wb:&\,�ͮ��k��$՛#�BEhn:���-���U���3��۰��ΪOr��H�6�70�,ٍ51��԰�A0YI
|
��K`·�o�%�Ry;�,����$q�d܏��>o񙭃%1���e��R0\���{3�I�-TG_.}�K26oX$_?��Yۖa�2�ޟqh��e�n�YPr�/�G���/�^���!~g���$5F񔹼��1X[�F!�;I8x�#4�	jt�!Y���Nx�ǝG�������'��G��s���̓��\�3W�Ȍ�G{�:�����jC�p��Ċ��ʻ"��>
�X��\�U���|ո�{��2���ٱJ
"޳#V��Ɩ��lό�O�Z�X�:tܞ4�v��ƫ����J��ؚt�`Hv���"�!�������nu�O3H�u��k騦v��d�bژ�l������wq��j� S� �2��3�8�q6E�Xp<vOW]�m��oi4�]�~�,[��2|��{c�%tssb�q>��%(!�)�X�}�/.��HH�4Q�C�a�`&}1Z��6]���b=;5�.!����C�Z��:��������n5�~��o�<|w�8O��1�+'�2us�O��|[BZF��� ?��u��xh1��6�V��B��L8�=S>���h��������	������f����M���W����9w|͒�B�k�/��m�^6c�K@�Z8���8B�tI�d����%��$:M��e������vU��s0�G�[�z=9|�|0�d�+�'ph�X�&-R琨 |���Epgqjl�q��o0b1�u?ǹO��3K��B�ٮ�y/ Ə�U���h=(�,J�}����nL|��{�B>!�[;i��f�� �/�$�c��ӂ�zR�SR��~�4��||��!=���-��JU� ��)|��w������G ����0 z֎G_n�xI���ԣ`�ӷ��|+��(���rrc���i@�MʞW?@[TI�C#Z6x�{��e�����c����x����!��/aK曓s����?��I͹��i���
J�K0�s:J
� `��B��5��o'<yz�QG�I��0O~�Ѣ�q�t�J�����ykӃ�_�i�2t7���JF�(�z�WO�V�$ql��nyC���A�a�$��g�>6��{.�aL	_l\����-�Zo����wa��'k�T2̓?HS���)�����I����j
	.̎A(Hkl�.7��pD������ʿZf��&�:�pT��u�w�<�x�c�����Nk�'�OrL��i��ox0u��x�I����럑��F1��JTLWX�e*��P��H{�R@��/�8��'����B3I@�.�}F��E

�@Ʉ��+��4��ȰIհ�	2�̌��HI\~�@6�?�-�W-����&����������ڜH>��^��DXH�:�b�5e�2#{
�<��N�q
e�$$�P"$6� +��$��#�xԳI����ޠ�aD@���A�Ք=^B/�.�T���Ԃ^Lw9���,K�Ŭ��|�İ^��w#�L���&>�ak�|���#���t_����������S����Eb<R���q�Oԭ��-���N��Ǎ�_�*���`��f"�M��<�6��"��	| ,^K��w�I8�"�Q2Z[ .^���}v2��0v�jl�'��)&��?���;�GDQ���C�L�(�V�B���ݱ5k�<��3!><}��}�]�,t�:��:�5��x�b��@A_+N�oW�@��vK�n�Ng��K6��[?#�&���]lA�H�c�7�Ea�m���ǽ�Ǿ�Nx_�#���(`9�D|8q=�ylK�Ѧ,�
 �,?=�'�X�A��lDც�i�)|b<��W���`��`�ܕ��C	��l�Aw
���;�>E���j��*7�U���i��ۀ��-�(�h�&�0�5���>��g��wם:��gvB���:��dg��jP��1��� ��0���0/�̰���c�Xl1G�3�w��hQ�2��NK�	3�e~FQ*�[iM��/$*GQT�58⊭z�l�r��-E8�d�(��b�_pnJb B���IN�}���/�����&3U�(��N�m��CfU6����{\���CE0ai��G�����Ʌ�k����q/�w�GH�rs���~&�z$�X����l��`�wΰ��6+��K�E�'XD��c��Q���9`�����5�Ų<�V��X=)(��Ep�t]FG�[P��$�3��Oi�&bL4�txa�������zW��X�B��m�r~�zO<m�oe�.��T#�A����g�1"�L{.d�|$�l��#�1PF�[��L��C"���.Q�r�[�t�����Cx��H���y�!X��֝���c�}k�B� ӧ�T���%��ޖbUS����e�M�O���u@T�,j�����K���hj $�ՉY��U���!�\��O_�ރR/�,���L�>�t�zZm��f ��Vx��s��MZL��뀪�8��I���}D\5�{fGr�ҫ��S��!˪*��1�r�"�יKr�E�����f�����0��@�J���[:L,��$p�	�9}�'Y���Czfǲ�O��*���7|��z�8�Td1;i�9��AU� QL�V���(�fI���ޱ�gAe5(���;|X��a��Y�E��=��/VuH���ܪ�F�7?��d�x��j��T�!I:B�G�;eJ)���l��	0�3�[�?�Ly�ApOo��J�J�rP��X�]+�<GoƮk��������@<�w�#lة�9�(m�!�����\Vٗ��:���FC���<]3��`>2�h�P/65��~�t���D{5�`�}g�L��9�A����P��?d `l\>��,�k.P.'�b,P�/�8, I"F������&ӌ��4��#Zٹ-sE�����__ |�y��zQ˵<� �b���`�X˓rb�|��o�U�5��+���r�=������)?��員v��d�y��b�_���Э��0k9��s$��Zp9���ҫw��*��f~Y��������ȍ���ܛ��-�PP�0K,H�g���e�a d��Z�gT��D�*ߐ�㡈�Ao��PB"��0�Lv@~��RP6��yHB�U=l��Q��8'�weo�V�.C��]z!���y���8�e�� #���r1�ݩ��3����S��H���X4m0f�k�
e�\����
yD
dm3�ze)�jk�
ͩ�
�,�e��ۿ�YQY$>[:?*�'�����Z޹榮k�|%�ڄ��X���6��LJ ��YF��{{_�@��.���(7��
��GM0�z���FΆxY]S}��n��N_ݶ0��߮ ��l֤�m��cg� ���XfP)�Dy�U���6��b��+�,��TL���tP#�S�rz��#��/W�e�><,i��J𐽊�e��`CW��}�>H��%Y��r��Z+����ǨT8z�1�)%@]�4H>��?����m���}H�`Bq����Wc=2c%K��۪��H t�"e5�pr�N���c��>��(��q(���M�'e�j e�6_؜�Q�]ޗܮ�~���%n�	�j��k�Ia�g�ã9�,�=>���p6�3�_��Y�g*�����4˒9 ���Y���`B��&�&��C��0gn.� 	_��j[J0�2��e�K{�"��ܑ���(A�*�Y<}8

�c�q�'f���H�l��] ��i��1`�$}���2��"M"��j_��ZFˡ�=V�R�j�I�Q<
�k�1��7,�/!3_�X��*O}Uw�XE-�5��	5EG
�%u��u �<-��^��Ix0ZQ!0]� M ���|Ɣ�f0%d�x���&6����)$ױ���Q�߮mw���r�8Z",85�+@ը{�$���1Go?���D?Q���������.C��3c�J���0�*=�R��[v&҈#�����B�C�hď�Wٯ�SW���HX�Z�R�䱄ђ٤S�5�T	�����B�j{��5�@�y�q>��?Hn{SЍ���]�����$���H�*�N^bw�9�E6�X��XOZ�>4Rg[�2��rHSP�ݵv�:�R���)�l� ����&����h�N���)�#�Rz�Һ���"��mD-r�|��W���5�y��Q��Y�ނ��z�����_��D�}����&{�	<��{1��H�����q���ycFv	?� _o_o=I$q����0��6y둸�x"U��_�a�
+�!R~*���`�m@5���L�Xl5"�:�\�R�c����2�ehU��Q�ȋB֬������j!lP�O`�D�Y�=˸?wspU�_����z����<�XN@ҏI#~[�|��y�@b��H��t!3���͟�9\h���:���|#��0��|����h�����-U���"��\O󣇻p!BdĆZ�*_~�/Ts�d��9}���=1����m �����|x>q�`��$<�&��{�!�M?G�rL���M�yf9�(M�\�&}��1V�3m�ь!�O���%ejh3ɚ�K 2j��P�@�n�ĐÐr8u������IN�#U��[��K��Ɓ|�pM���7��gS�r�m�r=��<���:,��Sbd�1ػe-�7���mk�����7��L�yl���JQq�ro���̱��G������O��co
؁o�G�U[X�}0\���a�,�����duY|�+��~!y(8Scx�F`=�d2� �dMٛS �pKC�*D�<�6�\{f{מ����mD�[<��߈1��-�����e"��m����R�R�b�.�NK�D����	|�����Oj��K�9&�0aJ5��N*��;�N���)�Ӷ�\�W�e�w��g�������k@�3ٌ�u���Ԧ8�i`�z�ý(��Ʀ#�F2���ڡY�IX��p�B�ib����gX�ѭ
t2�k��{7C
��8�:�く�y�7�3��(%s�I;�] �@i2�]x�\f3M����^DxK�|�l!���l /�`��pc� O�vM�����)ϋL��l�a�T:Ò^@ԒZ�*�t_\���8F���i�Z�gTM�O�W�@"���_�Ы�3M���x��SF��b����h,΍�+sO%_8.$�������#q)B��݆�.��~Ac=뎜����ݬ�'@_4�r�F`2�)����Գ� ��z^] y��������X�Ev����ǉЁr��xY�U^�ɿ���V�jH��o7�6�G ���z��dE����y7l��o�!U��'}_�����P�r7�����\T��pYT-��/�R�c�����*�gր�s��o}�#&'~�����(mѤRO�'`�
d�6 -�?���X�H���/���S�o-~�P[4ox�g�PIi�cl.��Õ�mr�!uIV-˽2q��zWȴ���\��������|y�E�J�@V3G�_惑��Ē�x'σ�6�h)�O6���A�ݶ3E�����ٌ��KY>�V�6
|RT�j�+�DE�eg�0�a�.�(��I9]x���u,u(�&����m�D����C��7Z/�PH'��U�$C��z���b��w���HF=E��Ku��kb�d��@Z�Af������m���v|�Xe�w��d��_�װi����ؔG��Z\f�P�4rȚ�m0.�X��u��ͤ��l,WRݻI��@�A�d͘����5�=2�n��>�Z�1ٷ�iE�Ԇ��d �T�@���y3�mZ�f�,��/�tU��l���T�w!`�g�:��u�?��y�"�A��âE#o��L\�
�6��c��y���>���)#<������; ��uD��eg>!��Gi�QQ�Y�Ė�Yg�G���;{J�J�lh���vH�duK�v�gP�O��\ԅs��v���ޱ�㤨� �(+�h�`���'�d@���5I��k�����^`̃�)%���"��%)f�{��I-AѺ����`�����PF)]�q{O�;�8Y9K�2;��Q�2^��^��ru�i t�w$ �t!y7yJ��{�=�R���W���Ȫͫ�cri2�|����f�&n<�~���Ƿ�x
�,Ŝ��/$4����S6�wq\&s�`�ͧ��<NA����n��!��&������t&�ܧw��3�c��+�^d-�^Ͷ��/����D�VRE�aT�y��2�Cf�� ;gߔ��)ή@��lqʀDYLoh{w<��u�#���_�u��/Eh� �˫�+kgt�^<u��!9ً=�<��r/6m*��͞�]5��]�l,��6��k��mG	+�l�e��k�Ll �j6L��R��"��3������+�����َ��wX ��QW��~\ʭ�R��x'��Z���W��Y�t%Z�;�&����������jw�9�!6��p��Я����D�Ḋ6�Ѽ���>֮ӷ�Yg�Z�(����n�C��F"�&�1\���L��V#��fyY8\/G�\��vqsP�Aj�����w%5���r�Pg����D(5�7�hH��F"��E9�Z��$�x�P�+�(�����b��l���C��t�U_B��A��f�O��J�B"�F�D�=CsK�G��*I���B� q`&9^Q�싕�㥘�'?&"�#��C��CMZ&5�C��:TT6](���:d��k�~�5ǥ�8��eōC0S_7���cG�O���B���Ś��Q`cR�5l1	M�w��.t�����
 �xt��:U�O��h �GE��ھ���<ܑ�f���
�?;]л���Ǩ�� ��6�������
3&�6�8Uf|��`(�0�u���̱�muhʸH�@nQ�󸒁 �������p[ǔ��k����棦< 9m�@!#/���i�lTcy��[	�a�fp;K�F��j��n5�I�h�|�ʸh��A��7������A��F�m�"_f-E�W\��	i�?1c���h?�%�]
��ee\���Hhj�n.�=���S&���(�	�P\�G���w5H�H��@vʙ*���O�!��B�6� n������U,�%'�Ѿ��*ʬF̧BzK��9ή�sWd�A@���:����98�N���x�7�{�|8HNX<g��-\x%�r-����'���24�;+X�%dv�X$0J�r��Ĕ�^T��BzN��c��I-OWڊ���hzV�����˞�YeQ�+��o:�w��C})s���G`C��w?33_mg��eƮ-��w�P\o��K9���n�V�[d���� �� ���|)0�YI(/ײ� Ӱ�
����k-�Q--J�*s,1��i�NM)S4+�;�����D�⢒T(8(yy�6��bdc2׆�&3:�P��^�~�FtSL��:P!9̐��ݞMd��4�
�. �V���Ɔ?�J����[Ml�й��ЮK����j�j�Y�B.c[�z��S�4�{`M�k�s�`��"/Tp�e
���>�#b�_�����A�	��T h�|`_�����LF-�>+��/#��~d�$x�����t�#�;�^A����db!Fb�����y�!�I�A�p�W	gaV
��mQ 5���ao���F��}-�Ͼ3��ZEQN��(k��U����7Y:TfQ�?�i�%�n}�$��j�p�����+%ȟt��GUu����kl@a��j�S�+�QМ)e�J�1���H��nY�L���	H���W��h��.v�]��=P?�j�et�SG�履�/���U!^�R< 1O��>����x޻�fk�=�O��fרUx>
���Т���^�NQ��&�ô,���9h�ͩ~E�g����)*� �[��X<�U��;����Է� ES�ma	0r�2�����#��&�@��n��v`�4}�=aDQ�料��G�XL~��S��(D��r���_t�7���
���}׿ofr���ك;�nAx��'s���e��,�	`�
jM�����d��>����B���j	��[��/�rH�5� �N{.��4��P����%T�
�E_S*�%���Y��?N��/��Tq�=�[����a!{m`ҋ����ק�=�[�vͤ�]�)�K���3�����<����	]ҳZD0�s11�
���_����5Dn�v`�G��C��hO�+A�nG2io]��}�aԂ��O��/Қ�\��c ��:u��Gm+.傹�� �GO�,�K��k���Fx��,ȔG�-��ND���p�<�tp�3-�x�9sn����K�`"��w�l�]����9#��Z�R��tò��)�V����V�"� ��)�+��ዑ��R�F|K������y� C�AO�}\:��E.��]KNz�'�p��r�Ƣ�K��6�7�t�]�$q-����cc�zܖ8[Z=W��iaiCQ3y�����:t^p-������m�n�n���� �6���e�R��C	��@�0$�N���������ެQH$D86�@� 0���N���]0�	P�b�b\~C�^��6ȃ��6Sb��Qk,�1��O'f0���pt�i4��Q���.�`�����ޜ �{�<�Np.��*./u��xbMC�e���ۆ�f���6�{�A�����6
���K�c�ڬ��;	c��c�>q�Z�<��sXKD�+�|���J����I܅I�`��u�����&j{���!PgKb��yd�*��8m�����s� io�LY���*8��S��F X�����G	�WX(���h�B��M����=��ΊN\��4�I?M�#)��r�\�,k������I��=2Ɍ�ȼ�u�T-�.�g�Ł)���ꈒ�ͺ��z3	�*5 ;�(�!Lp�~�>a�4e�b��XI�ioݹ�QM.��6	Tuc��_�sѳ�gO�L�݉<D����F#�ey㎖����`Y�y���z��u�}q/�`R!����4��V��,3\���ҳufꃊl���Z�ה#Y�b|ju�Lim���+�t$���3gZyfq1��4->���Ҽ�B#�� ����O�!�c�g	���{����X]͞�.��m��i�̔Y�&��P���.�C�Z5�?�0�]�m����t���������0�
!����҅	dbD�Q$U�6|�t�1��u��7mV�3�/-�܇"�xmt�N�d��`������mV6DW>�ڀ4�;���Dr@R����| �`�xЩ`4�����P>�И�H}|�&zh��ｽ��/���`[��.a(���Nv"Ҵ���70�.�G�2]z5`��!�$r�(s�=��N��	��z̺z���F;�lq��ܰVz����#<O�T_��s,�E�Kq�x�����7T�V�Y�&:=Zkz '�K?��0��9��L�٨�B�=@����j/#�˃Ϫ\�e�kެ���	�ɼQ�q*i[�2yT�,з`���5��E`o%
���_�G�v����	M7S&���?@\k(Qr�
i�M�ք������Q>�X}��;��\w^�Jh�٠ƈW�8��D�,3����c5�/�S�t�n�����؃��.Z��0�n��L�d7�A��}��u;�[I������۹�Ew#�JY;%��o�&p=�Ŧ���<��E^ ��Cr7o'�b<j̭����=��B�����M�h��v5~���j��
�0�����Pl��/���$����K������A���ݑ.��ʡ���&Tz�׌�Z��_���V�U����m�ח���v����I���c��ĳl�e���E�+�[^ܟ��$/Y_��II)�a�ļw�v��z� *��W�/S���{�D�<��C�:��n������]�X>r|� ��,v�{��+��0��[�Y0O,0��#Ck��˦G�:����Z��~�%q�"�����t9���}M������VKr��
.%��)�h���hĢ^o�~Q%S��U$��������y�]w�OUronf�h���|�@��B$�L9r8k��9������+w��j�N.�j�"h�Ȩ�F��� 齀��)����K�70�9��/*�26�E���e
p��2Ձe�e��F���⫨Q$�|�`��3����oB6��Ζ��,�CNhV�|v��ۄm�E3������iK�~Q%ؐ��#�~m��;qi�[}I�|-��q�������UU�SxAݾ���Ǿ*��"�/ZӒ�̋��@n��$��ȹS���{ù�H�/�Y4����a�6MHړ��G��K�L���aqL�T�0ic���0����@G��=�"�cZ�TT���ǭ�V�-����%C6L��?w�*�>�C�wy �5�%bE�38ֳp��/r��:���#��P�z��2�Q�u����U�~M����OU���;���~A��t�[3��ȆL��g#�y�� J|�����mBS��&j9׋��t��1��ޒz���B�5l�+�Oꬡ��R5ـ#yW����3���a��F��j�_�ELd*�o|j(�_#�]�\�k<�[F3;�	�S���:Cˮ���R}�T��֘���*?�q��v��}ׂ�����8��.���I�X�$"����1������8c�^�]��5G�!wV��V�<�	�erKL��������	�܈��"�%A�9��mM#�����sǹ���$/z�s�^�ߔ��P���;��%�}FG~���1��H�ĉ�����V����F���4�.k �Y�� w��5�-��޸��@\��#��!+��#}+H�Z���QX_�|^����������b!��:4��a�01q���������u�������(0$0i5��zc��x��s:�%|)��2��H�ӷ�eı���r�%��:�����_����(}p� �]y74����0�tY�G2�h�H"��0	e�'��ϭ����d�� ���.��X����`�"8:����B�=T���kg���ɷ�
����0�|���@���L��Q���?�����'J���0�䲋��8}�������M�|e�`����t ��
���g�v��`]�G�Q���[1�x��V#�@�*1|���(��;�����ר��tJ�������uϢ)���fC������z4�"�X��������ܻ��f���O����H�5�|Xp��HBң�������`���`h��3 ?w�	�����:���":��X�H4)e8���Ln�.U5�n�}�x��Yd�d?�j(6��J�?�~n���0~��=kKwu�{���x�A�ŝ=�l�1�&o1}p��6����N�U�kr�yx��aq��@j,^�`��o}ܹ��v'��Dce�pc^�my��~�%αR�U$��D�T��#GC��fZ���Jȝ��*��O�Fvd�ٽ0 �탁V����1��̟����4���^�֗�xQ@6�1J��9���!$�%1`6#��,L���*��Cw������U��A�p�C�"�����d���/���k|���~��i0�d!��L������T���&p�ױ�m2cx8�����{���ҭ�܋j�#ݖ��!`i���H,'�mI猺̴�If\jl+��<��z���7����R��;����N���VXM�)��)@�$��(���R1��B���x���[�i�}�%�`�c�����^3�`6p6�u'
L	��q\%б�}4��a���Pf����Y���ը�4��$�f�ϸ�l�r��QmB�>rǫ:��bg�A�^��lS]�>�H$�M��B�n5�\����O>ʌ.��04R!n�6"����ܐ�\�	2���tǶVh�[�]��I����i��v-M�V���t�Z�l]PK�A��(���y�֭��-8*�"!2��a��8(P4l�;���N���E��kxЫ��l6>YK��-�w�d�.�0�`�yv	o�;*Jp@�)��)A�0E ���E�S�x�  >��tp.� N����]��!����K��L������"�5�ey5��)~L"��_l����d������@!���A�>�j���D���%�n.���)3�L"T(prQGئ�{bF��9t�:��A��8�=)�Y	�2Vc��6\�%Ţ�QͲ�@��В�^y�F ��f���@UU'��A�&�g�d殛�sj���U�֕U������jNsls�n���K��b�����"�<̓�8��qB�jk�����2�?�9ޯ`�}sdF
�1�E�*rӯ��)������]9���� ���k�7��
6��]s�!��c�}���/�5:���BY�����!IB=�n��+���r4(r��>�Q���n�ͺ��>�S����~�}?��Q:
j<n��-��}�D�;����,��0ˤl2��f=�1�LI��²������X�@K���W�#2���8@@ީy�X�hW���Q�H�OlX(��iߘ�E_5�WSr����V$5Iy����{& O}�9��CI$l:��D�P��q�����dxwM�%��:Ͼd�;:O���XC<���0§�T��n2m�>ew������/=�+��������:R<N���G���^Pݡ���D�����a���ރ	��8��������t�������.S�.K<~F4G)D�Uw��k˳'��:|�@�ۙ�������	ũ���J�I����^5!`qu� ��=T�~��Ƥ�����x�/��S ׼=F��(��	�/��^
7SQoF�'�Q���h��m$X�O �K�� �[D?
��]v��	��!B�H���R�&YHc��E.���y�5�پ������ףi�FQ�e� ���zG1��02},\�#�� I23�M���Ql�!2cXA��C���JY�����2�Q�k��t��c��}�n�ņ��|)�djژ�ur�ٞ�RJ۷ }X͘��w3C ,�����i��tܹ2�6�	j������=h5N�~D�{�����.�����Q ��G8ayh1��V��د��}�\IJ$�ɀ�+���܅���e���h��$���%��I�`���M5?�2�	�s%���re���u�>�d�~?�� �nAY���#X����j�����I-�[H#Zx���_��t �������S1ǇE{�Ʀ�3��e��4���:B|�%)ܲ%��0WZzg��>��B��~�-K����=Q޴��mϾ�都�'b��Ƕ�t���Xج�IΑ�u��j�9�Cn���<�_V�q�s���Y��8����<O������|��0��)��A��b<���N�Uﱁ��ɌuTP#��Ȣ{�9��އˉ�/�*�9�v�44i)H���hX�8�r��m�3�G�WV���D^+Ubm���ϭ$wZu�(����}&'J�le�8���o!������j1�����|0Ne鱚X ������� ����t�5���L=v+�F�P�B�3����S��%�^�$1a�-���M
)��G%1M�O�5�es�rX��bX�KMw^ �O:�3��BP���;�HL(Q�l���ɺs:���ң.�G�LE!�S��'}Z����� l�SD)���>J!5����C���O�w���)�I;�8��`�%�_�(�P��ν�4��B���o�7�"��#��6��R]}$��_5�7���\��h�S�b.lB16��K��	�ӌ8:�o�ٹ�m��� �j��o��mv�.ph�c��_%f
Td>J����I�o�#-�Պ(c�_��L���þ����gk��b:/��s^�Y;\��8/0	��Xa|�ym�G��]`�	��D���9v��.����轆��P7���a� 6閃ewez����c�� ѨW7�[� ��9�5nݙ����Ϋ�!�X_C���?��٣�X1����-�C2!�ǇIA7�V��'��b��p���Ռ"����1)��o͟'$vO���������]6q&�d犢��Ά���z.d��%�$���H��'���H���6*�F>h�����>p� �ƺ�:�.�I�m�N7���h$�}��1�A�j�Mw�=��	LJ{h&O�܍�y��VU�U���Z�Z�VY������f�<2�P�H���Q�f���Ow�C�n�05����EK4{|SI����*Bj����'9��嗀�T���g�wSF�QFA��R��{�������ī��=���,���T�F�2]"�YID��?�,���o9��l�cF�v�9F�m����p3�{&�9��k���x��N��0�cTMj$٠M'd�f�X#�!'��m^m���Q���3��R,��G}�"`㲼ק�.B������0*[�Rl�w��Z�aU%шq��E]3�b�.&�<�c������/!3�J��3a*��(����s�$B)Y�����e:*�����a>qٰ׸#p����"Ɵ�1��h��\|g�t�wӬ��F��U�I�ǃ����tR�τ��¬	��>���7iY�7������p���rV���Z������o�v>7ɛ�t�k*)z�ړ���vV���+f�l^4F�l�j5i�)���.�rBfqm�&-��|]�Sm����]=�A��\(��'S�w�j6̱�|`ΰ�(*٨��e��
!݇Wx��J�fCW�>>��N�|�(�����|:\�fK��yV��0c�P[	��� ��t�X֓3AE�Fk��n �D��z�_��zz��JO:7�̰���z�1b����G@�o���cR��$��͵��M3Ot�-w�,#���?�/r��3js�zŭr��n'	.���h�YF��F�.�����:&�������5^$2DA��Y�n�	���@$>���ٙ/fx"�f��@����yͪA��q�*��9%�6x���:c���%�v�� Ǟ-X�r��������p�j�Ag���g1\�M{qB��R�2��<cc�cN���rDִ�z8��� ���-�:uU�P��B�#W!)����У��tn&n��~Y�=��ofk�k�P������;k�Z(�� �H��̄�(�l��>�H������C�@�oVlf7�\K�Q�Z@E�@'-)3A�	�W=f�m�k!��+ۭ�W+��ǽn��X��j^bx�3����6	⬿#�d��!�a��	���T�V��Գͼ�^��!:J��W��"9t� ����e�]�X�O P@԰�HF��9��&+�^��KlP�l1�A��;t�z�GU���E>�q��䗌e��;��M��ޑ���+Y�U�F����ϔ �9Eg������L��#�ϑ]� �J1�dUT.k���׉�h򚺕Ȁ�LPi�k��ڕ�k�ŇQ�܌ �M�-��=A'�rNƥ��].2EeBD���91��}�X���j�+�܅�R������h�}��RD�<J��2�:PϬ�nI8*�.�_���a�P[�q���7Q7��~�T9���dgG�tz�&gC�RЮ#�6��u1�M1_�.F��w,�Y�v�q=t�h�j�W��G�ES>�0O�m�/��=�^>8��Z�&o|ׯ]���#�����Y;�ԁԠ����_s�����#韽�_Kv�Vb�e0��n_Y)��p�R�����UER����LX�W�� ˿-��%hYP�7���k�<�v8�f�N�v&��R���R�
`�v��ʷL���!q��rъEh��EM]��K��5Zş����t��D�������,�n�;e/�#j��ś[Y)0x���q֤�ɕU��J�Mu�ܪJ@V��m��������;P96�E;1c��f���r�%A�_��i5�TX*v#�����$������E��c8"K��2��(��zC�;x1fc%����\�0���&��!��H(Y�����X�+�n��5������U�:B�{O�zo�iw��my}F�'�Õ6�H� ��fMU�Up]��{�K'��}��ϹX��Y�h0?�G�}���G,�yִ��M��-������T��smZ�9Y�+��˯,���@�К.u�O���x�(�ގ��
=�Im���TJ����Ƴ4��*#�n���*Qzm>S�'�uwe���Xw�G �����j��PJ-����������UtCQb�|����ɤ1")%�_	�	/yg#H	��(!�I��S7�=�D"�ɍ\��u�� y��$���f�JI���K������{�YFIGVr�� .Q��,r�+�������F�E!D��׽T��Ud6;�r�3v����&�8�r��(������=�T⫘���JU�؀�h$����z���	륀B~4xqͽ��S� ����9 	p����:���:����^��FY�I��!��+�OBo��Ug�пǥ�Q�'],�����=ŮC�t��a^�z�V�������[�����D(�9z	��C�=�ԇf5���b�ɮH.�P�E�tWK�>X��vQ�4�Ȣ��t8М�
�ܥ2�Vw�	6��:�9h,8���&]�D�6E���� 6vLk�ԧ�]�HӞ��Ի���f�7�Zj��o@�1�7��:
մ�5�괣��T���dk�{/����:v���Ԩ������`6n*#���g.P�0L��m/h ��0�.?>AV)��_g\0NB�Y���j�����8��+J���N{���W����+ypȆQ�T��
��:��������=�:~,(��Rq��"��@\ �^N6��`a���&�ٝ��Z�<>�ڥ!Z{��JoX��Cz�d�M�Ȏ�в=��� h���S� 9�z�6��}����c�A��p�ֿv��X}&�����=�'�<��s�h� ��Cp�I�4X��.a\��ʠI�z�*��7Xw6��Ԟc s(-aBΣi���Y7CU;6��,*�k�g���F���+��nS��J|���ҟ��_~� �������������j����'�ĳ)�Q�l 4��i��LM�����%4�E�?���Ǭ���ʰĝ�� ��6��j��6�������$y!ñAq�Z�C�k���|����N_��c��8I
�VQyu���!Bh@x��6wr��pʵ�Ƣ���;��$��:�w�2����+�U:\�l��\��`��}J�����Wؗ__ؒ�6<�����7�$�ků��ܔ��08`L���"����/$%'D8�=��KӾO�O*�*��i��+&��NI�Ba6����u�8}�ʛ�^����%*S�槽�P*��=^l"��E�5c��.E;rDI����U[�`Ϣ�j&Te
An������ߔG�/*�F�w�
�ʤ�gGQ�P��-g������������Gp���,^�X]М��ߔ�`[��Ǹ�w��N�1,����:3�c>�B�Q��(aW��p
�-F��i�G���z]�:�z�r�w5�4�s�a�̒���#�$u�*V�S��c�&a���QD�Ϊ���}��	P]�Y�J�Wby�&Ov>*���@��2�Lz{.8ᙲ{�(�$OZpj�
��e88[��Mw��C�7ׯ��b����-�����]
� [����+x��1�c�A�/�2Ѫ���
8b`hv�b�>��];��j�x��Ðv}����B�e�/P�@�M0+8W���{2�r]��3m'�*w�jꅭ���]��\�M��
nȽ�-J0����j=S�lM�B~�i�{Ѐ�;8��mm���SSY�v�d���j�'�3X�#>�󣔝=w�A�����d�סI����b�<��E�s'Y�ݕ�����F�����@+��T��	기Ai�
�C��D���>�,O�,x$�������8R-��U�K�.�%q�a��6N�aH�/\��㽔�����=tj�U�u;��	�ט�17PP�LJ��9ˆ*7)vtb6ǒ�T�ٲ��#�`,�� ���FS��G{0��0�i&pļ�r��B�M�@�G�)S�������u��sN�p��~��?34�G�\M���8_I�b�;�����dǮc�':��e�nC�[��hAU;�0s)'��
@_�Jlԥc�,wyn��W���w!(��%���~6��\�B���c*$�b���B��{6�� _���0���o��n���<��_ 	W�����g�E,:����oճZOw��JX��^QB�M��f9�KI�q���