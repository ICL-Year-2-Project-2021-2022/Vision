��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	q�v�Z��\R�w�0xtʎ5x5�������v�7\M�k���%n;c-<�<;�`.���B1�7���[�D�\�A��fIj�)����懋�f�7`_�%�E�i�j��yF���^�s�[wg`}vёp�M�=&d.�ȩ$7l	�$����>&R=�M� N=;5k�B���t��7�@>j�c�� �l��kyɌ�҂o�w?�x�)LD/@C [���"��ô��{ȶE}K){�mPuOF�<V�7���²�R�����7�?� k�V���Nq�f(.�;Z��)����1��}�mg#&_��Qo�A�"���FYč1+{k���'�eƽ ږ:���>d%��[ؿ���A��j�=ա�?dl�2�V�s祼_�
��$.�j�L-��S[l܉]Jȩ[��p���K/��N�OX�IE"5Ͽ��yMƅ�������9���:;����o��Yk��٩*N߰W���?�k��!��+T����|R˛�~����]h���9#�vN��۴��jf#GDPl��"�-tkDD��8��j��?U~hD[.$t����7 1��KdႫ���KW���r��Kխ��W���84"Q�2<��W�8�Jt�,�� .��Kc�g�8iS+>G����c��;;1HH+���j���ΈY9lܚ�4P(��!�9��(�,�;�q�=9C�B"�<���>�q��'�*HS�Tͽ��I� ��q0��4���������~�)K,��o��L���8@3�S�
���=b 5�ʹl<-I���;j\��K�(�wÙ#����#`Gp�-��Qn��ή�sC�n�Ұj���l2!���78	g��:&)꼤@����Հ`Ѥ��*fa��Ğh���U�"�Į�VZ���u��aXX̾�:h����Jv�y���^�o�N�X��r�52���kg�0��}>Tb�"��Ѹ���zɍ U�Ɔf�\���MS���TǓPZHРL$��/R1�j}�H����cKoſ�p�V\鿉�0��׫��ړe8;���ﵾE���mռ\	<a�;�N������k��!a���h?��y\1!���~x`��u��*�ȧي���$R��բU����/f7zB�$�M�%�`��"6�����J7�5
��a�S�I���a�J�&Y:�`�~ĻqEѾAC�*T�)�_S���@Q�2�v4�L��W6Q���.����j�9��&۠M�$e������}��e��CL�J�z����cg@\��H�ikۭgߜG,D?�d�Y�ZV�0��u%��yN-�	X��o��~��eb���%�Dl4
�o��
����Tܣ�eÇ����_G/Kç]�xe�maL)F�v斘��� V~���e���	��>�bz%�dj��H*'�K��� �3�x� �r�<�[R�idO2���"\����5�lF���o�׮�F��V^�A������ٍo:��aB��x�1�:��1�L!.ٽb����G�:SΈ�����v�h��j��gѻl!)B���$n�[��q0n/a���21��ARH,��˨M�(�`��R��WJ]_P���:�pm���E�T�P{W�n���^�E��%���	�uK�w���)g�fNa�;�"Z���כּA� 8�����)<�cU ���#�g��M�F�v�n�EU�=��02B%J�\���}f.��;geb�[���rG��O\\|e�¼pcx��b��mEX��]���m8Lۯz�$Ǒxo)�V�����:*��Ng�Ƭ^���%*�\C���0��o��an~s�tl+*4�7�;�ܡ:����Fu�D9�D-H��T�&{h�IptZ��J�d5������1��c�N�ƅZ�W�
^�~�CV�>Ql�!O+�#�;&.�ս�J,_lD-��NV�Ҧ�c��KE�8/Y"���p�_䵮�`a-x��M� #X��֛�V�@�))���Q�PG��4�oHvax�*�z�Gaon��w$���v��m��lw#���Y:����ӟ-�����H�;{G]��ci6
/�ċ��K����� ��|�#�T�U�'A������(�E��<��͉��u� vYm7^����9c�RN�
�>Ӳ˽<��������P�9
w}f�W��J���/����S��7�$�k�qώF��U�>c.B*X]yu�C�
�j@v��㝻�p%�;:�Sǽ?K��Ӿ����xD���~-_���l�k�rO�E#�Z�X��;����r퉀�]ZP�H�!	`�����Cj%�p��9ʭ�4�½�AcT�9/Q��p}bV;��(�c��3iě1�b��$)dCX��dm�ɪ���9�!��P�;���Q����Ī˼��y�C#Ͽ�;���[��fq��Q[��o���g�O�u�V�q�������(�jO�I��2T�@>�!ɡP�s�,���b�a�����V)H��#�T�fؘ�ȗ�Č�uٮ�([��6^�|i���8v��'��f$���^�~��?�'7L��p��~�����'��+7��5��	�Ĥ-�.���b!-��g�L������J�PA�U���c��޹���IS	3���z��@�!��c��Q����g��^˛���&����ԵL7R������mf�9�4��(@2f�^�f:7@����F�,$����4�ROZ��`4���f�=i�/憞u�4 O[�a,�7W!�-��x0�q�6���Dblϋ��p���|
6����d���,��ȏ{�&�E��[pT�R�Rj-�R�(��$��.�{{���NB�/ѱ,��7����6�U�`%ŏ}���w�����_d�7@c��3Yj��a<s6&~_�Ť�Ъ;�n�J�����ֶ��$¡�cz���<0�ͽ!��l�r��X�oWE�r+�m������G��I�ɂor�HF�Ù���6��8,�0E9n;LMV߇��������o�H�V�f{Å&e(�LCj9�P�Q!�I�aOw���נ�1��4쌞C/8�IJ��R�g��H�݊Y2Ǎ� �y��`ݔ&Цy0��K�Oq���_@���O �@f��2��2z��W�w�m�VG/N��X��}O{�^3�m�.�M� V3yų�I�mE��*�RM��J�Y��=ŏ�4�園�܃ÌVR?�L�_f0Gvpn�-)���MV���@�?Kc���pض������MQ��/=[U���h��Hک��{�G2�=�F2��)�up���'K���������?u��&䱬�_gg���*&��	�'�&��
ptd�xm `ޅ)J{	+�f�"_㐤P-ڣ���+��l�]��Xb�	Tz.�E���X�?8z:���ۡ�C��ւ�ָW�v*�|�<���?}W��x�Gq���ݴ.[R`��/����JD�>�_o��}S�"!���������<'���Ɍ�i�����;�I,�U�����j�?�܆QV�����us��p(NЁ�3F�F`�U���F ��˙SI����G	��\3�� 8�����9���a��P�89�L��3B���0P�.{(��Dk�S�W��H�3��N���sRg�Ng�틈fh�2+|�t�&�v�~<����Ԁ�.Ɣ�:��X�˹=绔�l���)bS�$�K������Jڠ[1��˴K��%9�����J	���Nį�_[xw{�W;�}�74��u�.�dm0�f�N�tK��2@��A��b�f�dK`�.�O�o�`�赕l�M��Y��HA�[���ͩ�p�F�T%k^��Ñ.�Ձh�#�cB�ŖO��eh��7��O�/<@���OQT�Х*d��+ޘ�{,8��jt�]@������`�_;B�X���	���"��Q�������R�{7�Bfu.H:"C�p�gg���h�-U�j&M�zT�"��I�����Ɋd�^�x�˝�Ct��Psi�aV��U�#A��ͯ���l1��]�ۣh��m��I>^�n[��9���ۘ��1�������{�sdӂ)�*��b�1-�&7�R��_��ࢲ��ǌz��tC�����v�C�1Q4GI:�FA7J��Pžm�VZ�$-��v���=$�{M�3O��R׎7�����p����q,O�@5��� �'��jx�9GB�� �����X�y�?K���Ǹ�E/?1)�����̓H���05�����k�v�B��|M9.�S��rW��ֹ��@�rO���i�frz��]8b���:	�U ��x4�;6�|j��ܳ��QGP�����ǹ���`'ݬ:�Ys�:�5f ��+�:�Ƈɷ��7����.QF?��3Q�}�9ꅩ��w���fv!?����`����Rm�߂��~b�O"��!S�,�(�|+� �sf�B�Gg��'�~;�O�/�cn3vIJ���c����7X�_\
}Lndڨ�u���S�٦h�$vWD�BQ�;�����C䞴q�tP�"'E" �y&J&��\�N�h�K���e�G��s�N���K6���X~�7�β����C"�I��J�mEmM`�L,-._]�m��5�''J�_��4���V;rS�9�Tg����{G�=�R�����������_��@�3��c���tV=O�)�Z�xVW,�A�mn�*�[쉭r�u�V���7��=�
��`�����rXM�b
��b�'�ZВg��-8�g� 	��@�22��B%���ޣ��'��)=�&�EA4�}^<H»I����م�ٔ(�ͼ�f{`<g��z0���:k���w����CV��m���E�yaQ�@��I2Q��d���4a�a����q�[i�6���@0�]�w	��҅�Pϙ��=�+B�˒m#�����KjU��r�i���)��J�
k.J���PE��# %�	D? 
���rk�w�->�Z�CRk��m�������}�H0�T�
�5����]#R�MZ|�8|�z(�W#����ecW�'��G��s��i�>Y ��(���E6�Z�� `!�C>ηcVbaK����%3bm��a��a�h�Q5�zs��̄�k)�#�<pZ�.3o� ��J�	s3~��[$�(U:ӱǿ�*��I�
�p�#;�B*�a
t� ��X�M!��}�����R0���E�ulZ7e0-��}rg��,�����2�f;ٳ�H.�mrS�/�"r�F�}}-����	�T���=1�v�w��Z��׼�\jQ���E1����5
H�� �ba��s>f��������3�̤2;C�H��d��AɑXv���V;���״�+��^^�������)~����������N��׍1��� ����H�&	�~4ڐy��J���s6�*���7B�!l����/[Te�E�mB�NZU��TES�ʫ��zm�W;��>d*#%~ǵf].�~�=8��Q��&�hN�&�w2nb�H��=J�׽�2�ƈ��9��)�zԒduf��5�����A�XH��W�/��o�!
��;�:�1�e<8�a`�$��7�``��]�.�<O�J�$!��t�qR�GW�C܃D�E��?E,��]�Ԁ��x����o��ɺ�Ț��h!QQj�H��Q�z�9cY�T7�Uo��c	�n�'�Ҕ�b�]�H��?� )J��5%!@n^#0�#�U��h̃}�7�z�#h���,�
�۴O�F���ii�u�{�Cr.r��6�� J�BmA쒥)w�ˋ�Z�5�G����̧�C�y#_*Eh���-�j�F_�%ѳ�@��3)�?I$�q��n}mt��oη	����۝�Z���G��Q�B�ج��bc�r���\;(A3�*{���!�;w�K���A�����4|���,G�^Z�%��D.BU����^�wG���ݽŌ�J�R�.\�22A��Q8�'�C�Ԓ�D����E�Y����S{x��"2XE�s�]�j�w''��q�-�H2pW����it[�d06���G�8�y�B���҃����Ӆ��Gڻi-)��^�0����U�l}S�ſxA�`~��A�x5�=Q�5t �����_�!oב�"�7�»h�|�И�Ve_�`��i Vἄ����`��-��S�z
D&��'����6qX���oķ�p�7u��l��W���$5�1ͼt�VLN��4��KC��O#��Zdn�񰖆��Y��!���拥A�n~^nʓ��,����R�}����$/[G�k;#uR�&�l�{z�� e���SU^�:��v��8�8Xjֶ�~��&�W�oT�/���}�}��t�kv�[�g�z4!��\������v�Bj�Eκ4��e������W�g�}�X�Dt/w �oA1���`f�>�(��3.�No�li#g]-?t!ehJ��J3]���"ܹ�(2hWv�b�
z�a�%
��s3Bc�(���E���q-X_��z�I�9Zp�|���*�ґ����-ڲ��p�<�t�3�E� �*��W���J����܉���ɀ9� 
�$	�f� �Or����2�[$��|4�J��%��0�������;ew�{"NSv�����׏�)*��?���� g��U����o�9�0גT�hfX���g�ǣ�\��UC 㷵�_v9���;���9���eo��o� I]S`D���\������LW�wt������I� ��C��=��7�����g������Y�)𽻵"�U��؁&�h�*�����E�k�+�!rSǜ��w݄J���0��� ����y�d��(w���/��X�DY���� ��R�e,��HT��c(��U����y��+�g#�	��n�?�(�٨���M��\��u�0���`t(l��["c�B4 Cb��ߟ�:
�+���d�r{]�)Fk��_H)��VnƵT+�Nb��H��^r��P�6_���8n~.�G��l�y��x�k�[C�<��ff1R�E�6b�禛-ܩD��j�����{rj����7d�H���a<�RV�XO7n�Ӷj�"�Is*zԿ�������yÍ����G���変X��̧]�k�\�^�m\L�P�o�Մ{�MLlg_�����9���z���E������p�3�]����Q�V��I��
r5���#C������-������h>e9�����[b�9��#Gi�
&=R�t�� �T�^&�F��3W�МS&Nte�s�I���0�i/rnG�[�ZYU��IR��j4��ȯ����J~��8��y�o�e�c����w U���ČCݳګ)a�\}B�U�>߉`6�����x1j���f"��$��;?J�� ��l�fm��0ܳ7.@`, ����8%�	�a)8�詹��'���{���΃�X=�)�7�w�X���	1�QA���s�9�"���	���]� kG�Zu+|���v��">�Mi�[@��N�<�M=ژ��eԞuJ�-�v#��8�gѽں/���: �ˀ�X��/r��U+��AV:��-����3��M��S�A6�$��6������Gi�^^S�wr��a+L�9�2�c)Θ*�]�:����/Y,g�ٳ����O�����v&�4�v���>��l�i�)k�b�K�޶��|�ԋ":�Tߠ�6D���>��x��ɠD|�aӄ�g|�k�ݍ�3U��.��j�d)W:�g�F�C�g��RN� ��J`�)V���:����y��J�k�	��)��sR9�+���1�x�a�j]��r�f�Y�eG����	q�����e�`��	�Z//d�ث�[<`��Z?5���H`�[�j���D���Z�ArVl2)
��>�u������C�@SD$��[�
yr���ǣ~����'рn/s�|h���8�;k+D#���!��@�q�-}��e��!LWCҗ51/��cO���i��Z��5A�͇��|�Oi�%ϛRE���l0�u�8�I�..��K\�E�vD�pD�5�2�'U]��*��uTu��[�R�+��X���g�wA�P����m`���wq��o#����U��E=XL��<�VidPP!�ńa�e�
n�ۅ�r�D/�9.�AM�V���߂c���~9����H,�}J�Y�l�'�EK��/``f+����4O��ӡUK>�vgQ�12�\3�ƭ�+�W ����V��V>f��g���3�q�p���?�cn�s�����'�Of�p]�(��������g(+ǎqf~"
� e[�v�Mµh���Y�L������@Q��/�~͉B�4��A_�X�<����W�*��L!�|���5@�7I���`�G�{�K��{<(�.4��y���Ԟ%uIO�q��P@�R)�NPl��of@Fͼ=Kɴ��&�Y;��8��H���岶�{Q�ʒlm��k��l�.6�<,8��V��@!��֥�lu������4~u{f�+�5�?���)>��_��|�w�t_7-�H��ͻoZ� .�U:.Y����4�FQ�fU���J���Pq���T۸���A$�)��JI5Fθǅ;�1�p�Gޤ{�e��I	c�����Ɠb�,���6?�Cm R����Wa"ߠ$%��q�e`����Z2.庲iL��ON��DN�5�-u���+��hB�Xv6��w'����Ѵ�=.R�# �l��w�ħ,s\W��ќ��רl��J�A�-`+�=�}�֒�03�e��"��z�i��x�e�9`�g�
� �*�E�ӱb�����
���G+��ǉ>��U�ŉ	59n�f���>h­V1�e��vIΞ�)֮�&��;��"�ۺ2A��l���Md<7{;�^1R_���}���W�K��|  �������5F�&���X"��\@�p�o!HkwɏK� �b-䎚W���Zj:�����Mѝ�
BA���o�Ȍ�u/��S�a���fZ1�O�&�K�&��x���6���;�SIź��ݘ%;ۙ.�!�\����Y�D�A'j>��	��A���AFO~i/��x5=1��36C����̈́a��d]2�'��Z�!�bg����y��7�G|���U��G']�t,th�h��<䑌j(���|dY���cD{O�6S�A�&M�s�B��>)=�� #�����:�zR�D�g�ٰ}iM����������߇v�>�I�z%K�#��T�!�.fN��LV�)&n��F�,w��鯊�mޡ��q���l�լ^\A�聄_}��FN�\��2�����l����!^n:�3�0�_r����KZ�5�
8#��jL�r��Ba}��E�&������ށ\⑜�DX+v�������\���Z��y��F$�n�[g���Q)\�k���k``i�!���X�Y{N"O=W�T���F��cb��Z�}�F��q���;�\����-^_}2`��n$�8�B�Vk<4R7���.�D_8�
�,��1k99�`*b�ۚ��m��:�(�-�ZY��ӑ����z������M Rº�8=!�HNs̋�-W��D�z-�J���z�Mz��M/ض)�����BuX���bsP3�`r�[@�͔bUYm�S�����*�ʇa�v�TV�?�ԏzĦ,Q0��l�o����g�藕`D�Ѕ�fb�Иɑ���$��
5�o�9�b	֔�~���.�5�؈B6��E��n]���m��L�6��/�x�b�:q���>��E�Y���\��16��mJ1J�@=�x����mi��Xە}Y��6��1{��i�ͤ��'?�<�1R�K?�G/�������+�֓E	40�
u=��tx���t�t�뒶��7
)�l�ۅt_��죊��.Xd��0�c��}���c\z����{����GU�ϐ����88X��1�c�8*6J�%:�s"f�J�X7��-�A�l;&g�_oF7K
Y��z:�$Y2�IU1�mr�������е���$��}wC�5<�8]jA�+�[W� a�W�lLQ*35sa����~�F��/a��##��'Q���j�V���U�eFk�-U�4jZ�o(�կ\Qh���_4��W��m�g�m<�-���O\"#�l.&�9�4(���j�7x����mh�gsf�9�k�>�>�H�y� h�f����K���(�I��@���<�q�lA��#�.���+4��"�o��~�6*�"<v�u����&P����|d�rYh���Ր����2�)���QS�/Z*[�lp���Ǒ�T$��s����B�YW��������%I��_m#!
��rхvJz��ﴱ�挅�;x�����-�y�wGe��(i��4Zi@���Y�%�X�U^�n"_'�# ��W&+ن���9�����ܨTK�"��!��N*�&�ޤi���V��.���f
�l���<��e�߹1����*�#[L2���T�
|�s%�����������m��1L���US���>��i�%������	g�>v�v>ۦ���:K��D)"�Uy³סVGl�h+6_n.��z�6
�P�եó���P��Q�]��vL�E�����w�]�_���,)���o�t{L�	�L.Pnȉh)H½��aŰ�+S�.��I?\��"�65G�Z�ڬ~���u��U�ОAH6�dv�{i��9�-��]��RںY�5o�����v��C��LJ|Y���'W~8V�\K 0!@�Re4�3�=�4K����u���4�TQ�Čŏs����);oqHb�XLjw �\@D4�`^���^v��'ֲ����:�	�NZ���<�����l���T�2���1�_d�ǷȎgP!ɚ�	淀�|)�����@�)��Sޮ�4n��?�9@���V�T���,W3C�����g<�,7V���(J���s.���P�H�_\�@=�%�]�#C��mC}lg�[�w�6
Om<en\T��:��x�ŷl��#��BO7%	1��P7��/���Y8�Z�q���v�.a���?:�#�``����R��q�u3ʤК9��1.<롂Z+��;2�@Pݻ+%,�&C2�}龜�	�����dw��z">�W��Jh���/���$%�I��){�1uP���zt�P�ɞ�i���
���0k�;����I��T������_R�VٕM��)�Q�7}db�`�����	Fv!Z.3��u�3�XX���A�s4�/��eq���V@t� ��1����x����d�3�vS��f>U��B��'�O0���f��v���[ោ���j}�fG䁆�?�T#�� �#�Tg�3D Κx��
\��;�G�u�a��y8¬-\��A�����ڋ�f�쎦`6� ����2���t,gH�>�o��I��V��;$YaWiS�_Cs0�-U��7�o��Z�l�	t-���D�!�&c����~���N��׼4�xH�Y���v�"�v�sesLr�9��h��=:�s���>��cȮ�L)�`���j�ɖ�F�[7Z*���@�u�'��I^R@���Fs�-D2�������f�zg�a:za�`��|u�A�����w&��sb^���tO^��=)n�]x<�nM߁�,��D�*}�]����`�w�@	7c�����sd�'�f9	(V��[��
�+k���'�G����M}vԥ�:̎H#�3����X�}��U�I�DGvg���l���i�6��5`B>�*EY֓������8.7%N��=�o�qu��7|�� ������;`�ع��<�ئۦ��qjg6Ӊ�@W��(�@�-v ��L�A/�̏�a�!���~ŀ��B"�P��|ׁ"�'���̌�2�"3�d?�#��r��R�Q`���@�Nz��6Nf�VfCe�ė�2�?y4�@p��9p��C�ؾ�����,�ϩƈ�T?��M�����5����^��m�޾B�֏<@�
F�BR4�P�m����Rt�����4:0�
��2zzC��C|���#ɺ�WE�FRhr����i�a�6_�i4�vk3?��rLR3�A��	�0��f���S�M�,�m�jzj2���c���ݳ�vݳ
yd9�O���������WTO�V/q���#��HV���m	������ڢ�=$2%�Ge@qu��ݕ�[0R�~�ɛ�bC
��<������9á�aE�V�K�	�����.Q����kn�>��,1�mH��J���ThiX�R/��z�ބ�3����`��z�k�YĒ���cTl�)����w>/K�C�G�,��1�?�Z��بC0�о�R��A;)7U�����,)��]|#Xՙ_�D$����U�N�5��\^>���l0�����C�I�K��:���f'����r��P8`��Gd�Zn�"�uVNl`/�]7l)�Z(AI��'�����2�N8�I�X_��Zm�~������*旻m�%=�D |�U��3dJ»�Z'J\�HC���]�ۉ
�O>�g9��aD�O���yT÷�� J�h�Eg�(Rp-��?Ӏ�מ8�΍��V%�My����84�k�9�yX�Y]��_�H:m�Uuc/�,�=�z�h˚1:G�����j�2�ٙ�%�$�����UNqX)�~�7m�����ϯ��<�{��ֽ��Ƀz��ܐ��;{�n1����v4�x�f%�FG;�����b-q����9��a�q6�&�o��D~Ed0�V���72�ӱpT��v-b��������B�K�{Q@�jAbx� �I�~=4�5*�ŋpu2i���2�����-�'�.�gXrk��n����]�Ĝ�=p:����v�
�����}���1�7r��e�-�%�ˌ+�0����p�m����%.7��!7��JG��ƌ������j��Un]��/ҁT�����VC �f;��I��x�^}�%x]�9n:��j�)���5)�+����"���
�h��d���� �|:�K�Tž�P;����g5/�+�	b�dkEa٠'!���L<#W��V�Ee�� K��+�\��E��C�f�-"�h�N�68z���U�'C����xq=$&.e���A7�-�8�P� ��-�B%���T���� ��̩>��R�]�x�K��!��+TMpLҐ��CH�"��f,Fe�>�-���`��侢���FV`���~�Xt��/���^5�8�ڵ\��z�m2� .���	%� a�:NI�� O<9f�N�6:�~�Rfw�1��pXLԬ�|�
���~}ܯ\P�z�A�%���Jf�R�Z*��Ȟ�R�Jw�a�Os��&��~�N}1��.����=Y�����:W�$���'��s�`)���?��L�L��(�,����A��1 V;2�#Cf�u����?�6R���.L녤��$qױ��/�,T�v�W����x-�͐Elzhl���Z*��[Sekv�����ks�&�7��t?]�X�ŠnB �� |-Ild��2��L���I��a(��М*c�EU�7fKk���	�e���M'�Um��\�+3��ʥr@���p�}�o�L�N��}�df��M�U	�J�������b����E��Mtn|I�$��Kˋ�Q-���C�z�`�_^������&ev�Vk�@<}�2������Ps���X[���F����@~eSJ���R'��u��CV�F�����
��O�	���,9�ez�d:﬜٥�.��ɏ�,�����~��`��E�Ыv�q�jy��b��s����!��꽹x
8r���z�T�?��5�j�v9�:�� s�T���NÀ�Qk:Cڅ����J�ٗ���^�uvc��:�\Ԡ��F��I'ov��	�����:��>c�_�˙�:z^�J������و�V�͘FJT�H����%��^����l��7:�Ĺ��� �����������Dq=q;���6���
X�IV�V���8�V�K��2U=H�����/�6��+��~!��9]9ǒ�����������6�ceu؉	�Y�)i�k�x~�:ΟNv�N"\���V�5�H�"�4ءx��
L1��`*h�X��{-b��W����t�l��-�PI�܈Np�&�-�7]'Y&P�ى�ϨK,d�F�[x��+e��3���Ԫ�j�?��V��vA.p;m����OU4P��'p�h�d�~ūf0Z�NC�?B�Y^,�	C��"���]Nw�#��l�=RY��D,���5�l�O�jO<�/�w�ya�LZ;س{�1��7l�\�O�0�?����8�:͐~��H�k�//�ώa5߄A�A�Y�Fٰ����c3�À�/Y�%R��A���.�#a%�\�����}⺾?�ۏ{��bAJk(�H-b�M͕o;1#�̈U8fy��F�52)���&����g`JǤ��o���[W>
j
F~Ev=y�����kP,������p4����_��Ǭj7��p��k��WU�{��ym�wh�"���e�Sĥ�f�Lc ��U����9%�NW)�4��V"�&�K�>�fں��~�xGY��[�9�����Dw[!�&4�-a5�'�����ت���K�6|�QLg�K7��C,��T��K���8#A�D$GE�b�}~��.iS�ľ��ۗ�MtT�ո�(6��)����H溤�S ���S�3�G���Ɋ:5~�gYR�Xo*d��-��S�D�8��F��.�5��u2��6Y��-V����a��E	Rj��U�����6#��S6����J��CTF��l4(���Z�%{������w6hz���g�Ц���'�G�P�T:K�W��W=Jf���%����,��̔�sk#:z:/�(�S�2--�@.Ybhޒ�v�_���s�e�u�a^joL�`�tyv��>�x.��udJt���ڪ��;`%�KS_��
��΀�?���J[|�����Kp��R�p��s��9r�	���N-hV����ё1������
*/�u��ې��_Ü�P�E��Aq�W٪��dc֝�R����iH�	dz���T.&j��^�ҫ�%�rP<�zT�^�S.��;ۓ-Z���20���XÛ^qC����'���
B�ÃeG�}�Ix���89���܄3���l��L�@x�o�(=%�����e9oq�Ӻ£#�y�s͹T��ib|oߜ���&�O]����d��@�b��� ��W콝���
� ���?fӰM+�u:�$�}K>Af�Ɔ�%���ƁK��(_�^/�c�����"|����S���O;�:o?��aغ�9"&ơ�r\��Xw�d�׆��b��NL�U!B2i��2�zu�lߊ:p�_���mc�S��ӭ�<='�()����1��i��L�f���El#'R�ޝ�XL������^ح�$ޣghHc� �=$�m����������i[�V٣�bf�<-߆'�����HDg�/д�� ׺�p;��?ާ�����������>\z���|��F�Ɗ|����JnT�,U�fA�x(S��Y��-A��M���	�+©ᆃ|��ȧQ�Ro��/}5
io��i�ب#l]�D�#M���B�^f�[��&�l�$��-\�3S��ص!�����	@^;���6�C�E��Eg���L����#�5{�W����r���|��=���LC�c��Z���ô�TB�06��1���H����ڎj��ܸ[�C�����c����SK �q���-�F��l��xʤݱd{���-�%��K��Dh��If|��ݱf�A���Z���\K���S�K��]��Sŕ)Q+�[%��A���uj��iU͉���<M���?kp��F�����2���ȟRI�����r��e�T?җ辦H�f���U �� 3GI�z�j�(l#g�nUE`��ޟ�}xi��#rc��]�4UX�AP�;��6�L����lx+Lw˜.3���y�.wʮW>���ضc\.��G2a+��߀c�s3�i��K����A��C�*����=�c������ak!�i}�H�r�1�?�KT��f���2E�$��C7D�o~������g[�C�X�ļY����ԩp�EY��v� � �h�Ȧ�D��t��EX}�SA�K�DX��uf5���~�x�*�>�b��ۊ�7ƀ2�)����j��a�?�OcZ�� �F����s ��7�pWD �Wc>���B(��'��z�θ���]�<�mӶ���8�N�^�D�'XX+���y��Gb���Ɋ��"�YY���'�H�)h���F��g#c;�`n����ǻ{���˪�lV�UA�7W�Y�8�� �	˲F�b�G8i�����#t��p~�6\���JAj _�'|�o�����Ϸ'G��N��
ʲ��,�����8�����.g�@0r�OAQ��#����T�qޯ�r^��� �̡ğUx�?�M���\T=�?&j�����78�������x��%?����F!��EW#���U�G>����+y��}R\�$a|�qOmH��+��ע���h��x��T�y��_y�h�?-�� FSVs���K�<T�S�_@��ð�L�C΀�a����FG�p����7?�f�؉�;�Ґ�̍A���}�[m��.Au�D���
l�vQ݆����+���J�/�,O9�y;2�vz�I���x�
����ؠM+�ȠqgyG��u�#� ��pG��_(Ԟ�h5HM��X%x5_����|z(u��� ���KB��U���+�QI)�w���΁шt#�꿬���}L�=/y'�ڪ�ʺ�)\�-?��"��]�)Gx��ҥ{,h z٥7�A�үzD�Q*~���̄}�"S:���o�"~��W�y�4��B_����[�?w9��-,V� �u����
�'�C���#Eї������C�;�[ɮ���-�qd�ߒJ̤�?wtf�Aѓ/����
5[9ďs'B�K��T��q)S.Z�Ǳa à/3o�:���w��^��l�w�<�L����xY�u��q���r[��H���h�^Pr_pÝL�5X(Tw�~	�74�����Ae�V���2�i�� ��`_��������wB>e�L��O.���#��nV�1�${��
���1�r�_F&/�@Qt�5�6�T�j[	(AEa�,���6�O��7m�p�[��ڜI���	�8��$_�,]�YҴX6���a�[��|Ym���|�I(���l��]�2�����Ҍ���M��s��I���Q������rP�e���xM�Cҝzy�; 
G(��Ɠ�7�[B�]�ĩc������T~B��
p`sL�q"�_�űV�=����?�O�d�:MZe�>I;pI�b�AL�%R�ܱW��-L�E�ep�@�M��De�i¦���H7�P&�f�VI�U��yA2֧~0S��b�l��s�������zj�5�*���k�"ee��r��vN��EI�vQwf�t��	4|od{�9<M�o���죋M����N��"����$���:��a�c��f�f��H��>�O'��l�� �l������e���[R9U!��{����B7���K�c����Y�e`��>���Q��S�V~�D���Ff΋`�Y�x�(�U�TI�W z�O��617�c�ݛ��������#x�uxY�q�e���vYѾ~~C��X��*]Q�Kb�u��{uy�r����#@#�|���|`�/BVClQ�u��&]R��j����Q�|WU'�teBu��.�P�ՙ(��H���ً=]�N �#@v�uYB���gHr
i�پ2O��u��@*����o"湈��! ��1���:�5N9g�`��R�ϙ�gq����.�OTXۺz��?�0i#��U ����h�����L���LN�c����l�<� ~�*r���Q{����O"�^�K�}���a"o稼�\�z['��'�2��)�,�����
|����E�zu�7Ls;�&jش��:(�3 b�|�OgJ�3��Q�����ٻ�� 7��PR3�X�f[��#�.i�W
{+��X4*�kOB�zP%uw[c���3���+��ԝ�e��**FGh6��9Kd>�|���hO�'�69���&z��a�OX������k�hFg���޳ŧ��oN�+�,ľz4H)F	i6����$���P�V�f#
n���R㣺^��7��}�밭:��&��Ҁ�-ܓ��U�R�$'V"x�(!h�}��6��!wmϠ���{U*��9!`+���b�c/Z���x���K_w5w��χ!9��_����	I�rv�։�qG�"v*�#H�<�s��B��9r��&{���&�I.O�8�Zp��a)��p�K�l!1���qR�l��b��W\)~��>e���QBl�*Q�� z��ݖ}6KV�O�t��x^����^G���5�������9|ey{��..�V�H�&�f[��[��Y���+]�K[�1��������0�y����I�L��㢎�1o�J҂���54��fx	틓a�1Q�{��R jÿ6jo	�A�v�0ϕ]���K�xC۠`�"���''}���DO��:�n�_�i<�4�.4�c4�.t3F�}+�V��jz�y]�TӖ��.��8;G>�X}8���s9��}yZ<,SN��O���Ud��,t*k��7��S��;�t���-k��@�v�{�-h�8� �}T�_+�������*�8����iz|��J]��>-�<>������ly�8򢲰����u�x�m�s��z\ qИom�@9���q�ى<���eu���@�7x�`<�O'#���@W�驪+�
쭓Z�٨%��22�6�8�5���Bh�69G�
N����Ʉh��L��ۺ�8��=�V^	��ӫ<�w�d�Ex4������L��2�K��~�MI'���>9(a_E����LL��S&+��J��>���/�hz��_/G��f��?m5U��P�m�Ā��Q6A/,h�=�λa|�]�T�z΍�'>�;v�qq+�~�|�f茙J �i��C�cW��~3E���Ч��g%� ���@�5��J��.3#?@w$���Q���x!�z���������FW��G�J}Ԩ�TY����A��l�H7w����=�΍҈z��-Jd,/�l��^�g���[҂��L�C-YL�P�Δ�u����TOK�C�{P���s3L�M������I����:��ul���Bm���x��կS�N�f��
��eu��k&�����EC8�ʐ/�o	���e��($xemy�_)ڻv�s�V2�Ǭ���]KY�=�u�Km0�u䓭Nm��IN��'�4�{08DcpK����Q��NkT~���> -7��'��,����Zbq��*W��'�~�:Z�����.h���S��x)�6��9Q���%{DapUp�N����s��6�}#h@z�(h�	�!�ґz4��>L�=c**rW������������f��b���ұ���-s�JL��:�or�̲���}"�IE��m����9�0��ݾ�z�V��������t�b�op�lo�$U�����$�@V���0��%/N(�h��d�2�Q#��j��X�b��ێ��(���Y'`J_� (4�	=ۮ�b��[\�Hܕ����k�..�{S�ئ����c	~^hl�����6t��#)��<XXy���e���}J7bR���B�P{52GC%��I�4�����{��d�ⶱ���&ip��n$��;	�ݾ�6y ���%))0w#��n�uX'��L�&�0�<��:��.Ц�Bz�����
�����ţO*�G��J}�̿)�����E���^���_+�[y�0����o��<$�
7�1y��	̮7�?=�.yS$4w��6��D� ��nڇ"JcG��_����[~;%�"��.�SK �mڪΝ�0��ɯ'�f�E����ʀ�*��P}�P`�-�5��+��	�Z��<�cEBF"��.��+���X���|��}���^�{cy?�e����^�湀�
�Fɼ���J�>kS��A�E5�CU=�����t��=VB*@:�bz�Ot�V����ށ7�������PF��H�z)�
Խ�^.<ESL��"J�
�������GV�>���FQs�Dݏ��\��*����B�����e�
��?��RHC+��e?|X����
�fx�C��Y "A��%�7�p��K�� z+6
"{mhx��a������	�9h\�-N�L���������3ҡW]���{S<>�2�N��=��+2�A����emCv)]'�ݝ{x%+�{#�&g�|��~MC;Ue�`'��t1١e��30����76E�\z�DT�������L���w�H�?��P��&��muT�ҷJ���@��dv�ħ
��һH��wqQ�1�2�W�WY�M>�$�ܭ�=e�d�3:٢�5���k8��
�}��i�UQ@+A^�}�΢,pF�@�����IO�Ż:�HTQ �эҲC76��2λV�!9)��%Ч�:D��s�����4v�����s��n��S�l���G��3���ʜ��4vKy�:�s0�8�4b�0>��̈/ZkKb(�h�F3O{�pPmDH���1�+���>J��F��w��±d�$9�Do�/k ±c�2��$���sD{ƚ6P�� ��gx8�w�gq%����He�qOᢶޥhq7YE���ܑ��bЃ	�����u~F�c�`��]���8��m�	|���ob��8�����͂���(������R����1s��_�����v�um(�'~2&2�����)�z5`u��� �a�N�%����"uk��RJrv���ېI�vo&����(+�w4i��bP�������O�^��q}�����@��S��i�\!ys儨jQk\����x��H ����Ur���cc�]@���Q���ܘ�J�����$�1��e��`�p�0mL���Ab.��z�|��]��yw���I�1iV�"�#>:�J��hH{�3` ��"<��o���]7�IW-���!&|"�r�Jf( hj�s���]�>ז���h�|��z�UV H�^V�h\�9���?��9��u�+��W�u:{a%1[ ��b!6��@@�n�����P�3y6���=2.���[���r�w���:5���w�!w�˴�����[�:���E��X�a��w���c��'��ce�x>ԤF�)��Ө�xV�Gbu>��%v.Y�����	�� �P�Qwk�UodT������t�\�N�\�M��,��g$�Z���{`[��׫JS}��y��JT&i\�g#���i�z��
X=���0�Md�a'�P� Xd}hX��4P�X	l��W��t����Ê]^~>/'+����K4WE�*��#�f���\�t�ri���U������y)�4��:�O��\�R:8P�JPw�X�*�����5E�7�(�4��͉���6���L����(�����4ȧ�fŌ���'-<��.w��&: �ڙP`'�'u�xО�x���4l�f���
_�x�&&&�����jؘ ��L�y����|çK�8�v��qG�� ��_B���|��Z�B�v�|��y���ry���8�{��يd�Y�J��6M��\)1�J��
����͇�@ۺ*w���puP��/�T-���4D��iU�_ą���+��n�@y�Aj�J�b��-�9 �$�lu�O��h�^ÍK �w�[a]0
�Y|�W[P�,�jxQv��Zhn����m��K�P����D����^�?��s�&�vv�����z���$ۂ����
C��]ݵ���P@E�6�r�/�������9�Q�jU�����R+�;;�JG�X�DO=֌�n���c�oҙܢ��eM�V5�ʽǊJi6b����=&�HG�����F�J�tC�8j+�J8�V��IU�We�Z,����Bώ�"���u�M�����c�7p�x����.���:S�)�ۧs���ːF=�W�D�1�pB0�9l%Z����V��$
7+ǥ��7��u�~��F����j(�@�BaO��]�z|�v�2@����YؾA2ן'#��Zi.�������̹_�̿񮳢Ay���AZib�B~ĝ�W�� ���	�n�Fi���PM]'��7J�]ks����]-����'D�
~H��;�2G�(1(��%�u[{&��Ӡ��iV� E$�pU)e.����j��%�<>��WS��HB=�Y� $���{	[w$�!�(V�oW��G�k𪳵w(������z4��x� ~�a���pN�.i�G�׷������iX�զ�}����8$��_��!�%�N�Cf4�z�o�e��L�����4a ��	a/(��/w��(eC�Q/G 
D��G
2��@���L���d6�56��Q)g���G��A�&�Gor�W����R�|b�!K_��w9�0.�vy���:$���
�`)�c�DDR��H���|o��ƒ�}H�,����]��kZ	�)/  O�~O�#qƀ'�Ɯ3�v4�%;
T��w�(7lW�U�(M{�G+�lc���>=��4���-�Z����G᡿ne�	`ç��B�J���S޴W˵�j�Ïh`��+m�;�>ᦆ+�R�*~�mE1[���[�@8�K��3B	��C,����@*��6[�/j[�CU���ҟ�S��a΍yͯn�U��:��쾼��%E!����j���r� 	�9��u$�YT�eƅ�N@�/���hYqs�I������-n��`#�]2K���hJw����Sʖ���)]�Q�)���%j:D�Ƶ��ϕ���X�|v�X�pl��J�%��y�P/Va���gi���5k.�i��/x\�Ğ�ۄ�V�luY3��B@���эG�SԞV��w��TW�F���AV`�wvt&}��_by���o�~�ɸ��݇`[ʠE������p�gqNpp@+�|��;O9g�¨Ak��o�����6q~�R�+��`�jY�E�!���W/ӛ1`�TE �w�IR:��A: ��/)	)�.*�����BqLi�CM����U�%#�R��X "nԓ�P����]B�*��.Yg\�t~z�.n��eiJI�tN>�*�@�HIgY7���Y��󼜑�a�`\����B�v��R+ȕ��	�_��7=;�ϐ����v�9M�*q��rD"�n��@t��z���7yr�����\tH��[��S�0n��n(�+g�*E}9�p�����K]�C��̶R[U���91�t%��j��y����.:uX�J煾x���J�lP�%/[ȭ�\˓��h�<韞��� �������?.bQ�	)ȯ;�B���_�W*2;�q���٬ބ�z�N�}�>�������x0*F��2ޝ��3[pEb�vO��J,�1�(�Z��� I��Jc�=� ��\���4u�b�� �/��m��!��2��?]#�ŞS�f�ߑ���b4{� �nZ����buQu xa}/Y��=x�<����[�^�t<=<�<����3}��8g�|u���h���{+�r�*�x>��B�s���R��ri4D"r�O累}e4�<�d��0n6 :�T�1���21V���@N@׌A�i��O�U�C�O��&"Q>߂3����<�f.�sAE�qYv.q7 �����[���Wr;���M��lc��G�W�H{#h;�zV1��/��n|��Oxo1j屯�jM����Xgͪ��&���Yn����É�����Ҝ�V�-ru/��r't��p��rl����k��7��yc����/̉Y���֡��Ç�7�ǲ�/�W�g"�9�B��}�2��(��#�Y{9L*�#Ą�Ҷ:'pj$H�l}U}���?���ƼJ0�&�h�v�Nz���ùj ��l�bV�Tomì�����@�>)��p��j��V�����Y8�-CX'f[�{
j,n�C�%D�PY��~޳�z�w�-������D��� Ro���cPUOc:��c"2h*�z�2Z�g���-�O����Q �7r7[�K⦊9F!�d�v��^�jN3 5�����R�XT����i7��>�J�)�8n�/�u�9�̞��V�Z,-�F����A���w�� W��͓H��� 8�m�R��p�q���O�<P�� +6�V/���`�T����)Iz�c�1^�ŵ�>N��Թ�G/�L7VcsHP���Y>>F��V��
X3�g�yǶ��َ�*�vai�x)�q^ϐX���o��b?TZ�	�����%�K���v��i��7��8Y�
D������+�
N�~�e-�wz0�D4[��4�>�p�I�6pJ�����vb�h�K�w���5Jޡ�Da�vn���B3���÷�	��8X� ����'�3~n���<��ker����A�c"x��o�d�����9����ɴ���%�t��6��T�#�Y)�͜����`s�i��3�Თ�����Et����2{U���C��!~+(v~+���`��^�/��j@���Z��وڨϬ�=�	�l�o�]��+c��Й��RL�wjѩ2U�3A�`2��pO���bT ��1� s�S'#�R�S�� o8 $ F�Ql(T"J�*[�k�r������W�׊�(銆`�xk�# .�)���ˡ4�@ё�׎��Cȷc&���ع�n1�/h�lVc�D�xG�!�����c"=k�Kʀ���йŇ�p@���@"�k�b1[yC��jd�� �k�� oc�X��f�~1@�cK3?�~��@h���kQ~�nIP�V3��g. ��I��R	���� (Z�R9�X\�PT59�v/?�nu	#	~%��V�(]h��Օ��	8��Mj�#`�I�a]�n�Q�V��0�\*�44}(�m�v��9.n4bZ��L�g"y|���Zx�.��*��1o�W�\�� Ahp.�?���p�h��$YaO'��}�i��χ�j\dz��f�;ٍ����l'�o���s�3�X�=U�6?��?U���"�5:������_H3��0�Uq1��<�'���x��7�3�@2[�`%�Il��Lm7�K��.]5�xҵ⎂�2XuɃ�����0o�x�(r/ǅ�	�NU�c �!)�~��Bݛ�b/u]�KǏNY���靣c%#<���S�(y�����L�����t4i�(�FC��ٙ��l��@��Ur��j��W�M��T�Fڅ�������$��V\8t�y|D���u��m���*�E��J��
J�V� �&�����UR(a"�|�#�ǆ�o�jއ�-�'Rĭ�<!ͱ����ֆc%��.��hE藭ս���2�d0w�u��O�I�#�7��ƌ����mo�ԭ��i��RM��x��n��&)��At�~I��2�v�h(	�v-5��YȜ�VE��rӭ�-�7	c�����<��^�q�o��6.y������c"����$]4�8����,�}���
��+;Ԯq��$�n<1E���C�_{� ���K0b~�Jק�9;��Nqk���wn@V%��h��5�yh!y�ˬ�!-q�Ņ�w���I{�6�_-�nk����T��l|�ޱ�+��&}ӿ{��h���$cTʛf���s!$ۥr��>]+���ۂ���S��$m}	��b{,����eg�!+T�}��fmTܫ��
�t�:��#�IY�ۖ�&��z�����-��wX����/Bn�@:Y<~�|7�8�m;��˒�W	/��0����KK�FC ��dSh��,Ҝ��Q4۝��~����{qު'�{#��$Σ]���*�U5<����^?z�IUh��\3��Xh��3:���c _���J%*��%�s��{��݊,9�:?�.�$�XF�n���R��2�!��RD��Hڿ��2�Z��g��Q��VGp�z�Sɡ��њ7P4�s���]��QX�fգ���VZ8G\Z�}mN>���6L�c���SElMKpmg�Wxf@�Иҵ��$��R:[��W���Y���nJ��}Eٰq7[��Y����i�Z�LLciG^8�Dc�˼����Ͼ��N� f;l�E��,�wv\��T\Ty��-���jŹV=s�fc�x W��'�Qw ����8X��L��Th�
{	��^��3��+�R=���� �u�s3�$T1����k�d�6�\s�l�0��ؐ��Wx����̕ ����B$RJ��5*�F&��-�߈��e��ޡ\�y5�kz��i��Q�%���|U�����G��q���b�l�]P�AJ���x�N�Z0�K�s\�W8M
c�<�m~P,u��֔g`�-f��T
`�4�h ?�/tŉ�c�'����s�QΏk�w����"��� 4�^�� ԡ�;��h��~��:}����2/�Q�d-����㗊���<(�B�U�,Y�Ό� {s�� ;i���~/ ���촚�X)��9q%��~��������4�;��Wo��L�gB[�2��`FI�x�ؖ�D�yM��ƖDZ��#�v�{筑E�g�/x�*w����5�޴G'�i�Ũt;Q۔�T��ܟ���Bk���z��m��,(���������nT�9�!�V�A��aJӥ�C�e��K�
�Z���}��*u.��R_s�z�U�+F荏.�}����������;z��ٌ�^�k�� �=�x��c�Df�_��9ҼʆQ�v��$Z�;g�׊���/0��H��h @�y>%%�d�'���7z��ֈ���1r��D�[=n��8��L��G�jC��Tߎ�Cy�	�����K��o�?�f7R���Zp'FL�֪���o��!���#�@����\nL��ZAX�i��}��8�\I򼾌H�c���0�[t����G[� ��U�ֵI2�#{bB�p�Y�S�]�-Ҥ�ք��L�|B�m�-�q��x��ߟV�ׇ�=8K�m�-��T�)Ƨ]��n[��ȆTz�	�z�IA] l�Q�(�I
l"}R�CYf�:�Rt�m�ʳ�L�W�Iܻt�Hu��B�:����D�����KE[ʦ�1I��I*�U����.�����ag��]��A�Ƥ�KT����Ç�nxT���n$y���֫r�����%����j����X���m�!�u��q������*��5�5ek�_��? ����U$��V��h��̞$w�ud��"Tc����js�����J��ϻƤ�:��$Z����#�0�����уc�J���[ͯ�d��:Wr.F�k7��0�A��r�@P �Q�&�8ߕ����~0�	�TJ��MQiJ�N|��x޲nt��Y)3:���q.P����nu��[�ׅ�"Ŋ=�RK�3 �\��:��c���On\��	F���������D��L9($A�2��Fp�7����*�O�s������I@��D��!����vK�QwkQ�d���r��yg�H��z���L�oF���Ti:5�;�h2uF��W�<���!HM45��~^�2z�x�3û�4�.Fk�X���*��eݐl���&mw~V�!���+��+ -.�\�󆝃�����%�N�1j�h:}�Z�:��&��a:�o0>š���*�B�[m��a3Ǐ�*�KH{Q�J�72'�G�`�+] ��~�o���6�Pb��0���CP�q��&��}����@tL��%śP�{�a�j��u��lغS�J�v�w�'��J�	EP��x0��ʯ�7Q�hu���YGs�m� ���|����!l�����O>�O�ko�kJ����L)AXE��H��D�Ӑ1j�B�a�,.$ϻǖ����%��O�8F؂7��X0p#����ئbm�ac5�h�8�M<�:�%EH
�E�����ʓ�|�;��߹J�(�e�gB6 �l����+��"0l5���&�!�h*f�-�]@�Đ�~O����6'�Y�}�Z�	�9��[ԃj���K�!�:ը����?ٍ��擎��	� ��|�p�vH ��EX��X����6�7�^��R7T3R�H�����A�i���l���@�5uPZ�A';�-z4	�w5��Q���^�a(�x��!vǏ��_�ǝB�a �!�Mi-�S8�M�Y=���&�ۧ:="��$d����{��&&>F�3��>����Y"��QV=+�c���!šW	
M�Ù�~ay���A����2����\΄����O��w��/��&�֙�
��6���Cdv'�������lV �Gr���C�����ܣS�v��d\�a%�V(�_�G`��*f�����Н.�e0ġxAK-8�G	�W��c�N�mb[
���cj[��;H�rE�N�I@�^���N�����P�0MJqG��^�Tce�qhp
�s�?����rB��])�DSA��rc*1���v=/6�>�5�"�1$�m$�0���6�$m�����?�ʦ��[B�#:����Ən$߷Lj�=|�&�V?�H��)�H�"ӥ�z��R����.U�^�� %� �(��z��'���K�~���D� �zB�~,c�6��ؾ��Ֆ��o�?G�xń�I#�.�k|�!��Ѿ�n�������z�@����n�g�b4dBt�ߢ ����Ή�c-�;�@���iZԋ;�Zj(n!�$�7����wH�~|��*�ㅵ 14�v:J��v�5A:^�e�1)�(�&�g���s��I=��#[���l�V�+�
A�.+�aϫ��1'E��Ϭ�r_�#��ʕ�h8����>5A
A���Yށ�YOV%��Ū�Zۄ��J���=�wf ���AI��b��� 1������IM4-t
6�}ok,��p�Z��5].2`]9�>x%åV�yi�bo��g�+�:�%̆N�#7�^�[w�����_�t����w��0��5��Бt�u�G�� /Jѽ*�@C�l$��0g�,� �A#$�u��@� �r���D�-����,_��;ʋ��؆Y���d�y�蘔 W��ۥwe�hkQ�A�����H>�XF����nD[�?��|�Z�nH9�
\�>A�n0�ZF�N=�A�~���k���%O�2`���,3ɜ��Π���,څ�H~-���]<F��9�kCZ>����(Ĥz̋{JC�76�Q�a��XPg�6��'�!�������S@b'��ɡY�YSx{^ፄx�k_:�J~�MO�~z��j����$�&��m�ɨG�C��Y.( ��`���9F�����?�a\�&��|�����?i��wu������0\�@��
}��NJ�,�����z7OMA?���x%��W[���EW>��i7�Z��6��Szr�s����k2_HFLsc9�3���X���M*j�y�-܉ ����!��\X�O��bY��s��r}9�Z�v�҉
� O gʲ�z�C�M��Yg�n�]��?�eKcvLq&I٧ȓ�3v�����@ه�Z�G����[C����iQ�VΥ# ��n��r�.0@ ��|w�)<h��D�ʣ�m��~&`�'�,ot7Q6�Y���u���%�����~�0��[K3̀qh��V6=U˝0�*d�Fc�}��H27\�^6��!�f�>���[)dK���4*��n�,��IZ�M���xW)D%%[����o�1s��z��AI��I��l���z��+�4Th��MFH8����U{�۵=�J��4����UK�=	�ũҬ|ɕ�ۛ��@��笀;������;ޟo��2Z�k��P��'�HqI[�Pq��f��CÕ���d���&TR c�a��-���>a�"�	�N�k�5"��:#����P[��o�14:�O�uO����cɗ����	�]���V��_��?�Kޛ���+�/G�÷��S40.G���w����!ٖ�D ����x��M9��� �7�z�<l�C&#��ܳ%8;�z��i�#or�w*nE��&n8�6��kn���~c��n.���Y@�F�Eۍ4g�x֐:��U�[ɥ������pB�d��X�H'�R���i��3�C���)!*�I9����������<a��{i�}�����h�9E:˩)�=ɐ�!%��f��%�����9�FS��
������0��'L)-l���4��,ά�-N��2t���ǌ.��Z�Pz�`w�~�`��*A�q���RmߦO}���P��sk��Yҳ���:6��"�o�I��h��E�o�������ku�c��a�<a;������<ҹpSy��UT'�����W�����:f�6 �m�$u�WG���j4ʎR��x�3��9�J���y��T�%��_[�5�N�{�&����:R3�!�d��ĚY��au���,����] �
�ʧ�n��:���E�U%�Yd�vS��2��YE7�E�V]��,�ݕ�՟B���>ϩX����@$�"��U�nP&�B�}�+�
�^��h熵r�t.���n������t<�-�uӽu˓�%���V�DRI-�^�Wnh�9d?-!jby��3fKбH��M*���}�ܘ��NW��Le}�:RK��I���} b���i�2�p�"b��hTR��P
���������Ճ��1�d_��me�3���f��0v��v�{��Bzye�-[x������.c���������#Z����s
=
��-�E���Q[)��K�Y�5a
��i��GL�/�>�ZphrXL���AP5�٥��z)/e��8�
ܽ��H'1�"��1w0�����e��1��}�1&��[�����B�\�ex~�UԃӨW�(@Ü\G�Jl�Bs80��zh��	���	�1����7f���I�g|	���+0G���X}�3��=��y�tdق0%w�� �8��f�T@�����4&<��#_lK|��c�nS��U(����K�`/��tX��vZ�X)�$h�u��$β�(4�w�y�7�l���ɧc�	Gh��o[���b7�O��C?��S3U�Ê�yWa�����[H>�~�Rm�`,�1q���ߑ`kء�/�{㲭̅�?��Y^����a5����ؓ�������*�~�;ā1�����Č�$���C�t��܄1�O]�o�
��^�D6z]���P�<�}�ɬ�ަ�N��;OaaG����"_�Zt�-�6�La������co��pqzT� C! 2�	(bK֋�l�a�	���:�ٜ�����6-�!���]7�0j},2��+�>5�X�}Y3�yN�8�4�ͿO���Av1� �5��s�4\>3Kcπ����BA=_����Cnw���<9כwL���z��%3�f͸kK I�?��T�I ���V~�Zy_��u#���զ�~���x%��5C�L?P���y 8nh�����ۏ�����`�e5�6Xc���ן;�O�������X�M�=����E􏶏����u4���K�q�s��*�X���p� {D	
�6��0�K�U,A۝2���b #H1���/� �y�̑�����^�ˎ ��Vm:� ����&����m5����ElNdj��j �L��6P��}���'�9�X+U��&&��%	�n�M�j&�a��p#~t�fp]rM�=w�`*��J��t�<H?s�V��t�1��ք��x�*0�Jש����Z�:˾=LU�U�5u�$�T	��^`��-AWY�m|��1���,�[YU���.j/9� ���*G����_v~O�b��?J�a���[|�	�Q���<���T単p�����1�9gxw��*��l��&Eno�W�\�1��;�V?�������]6Q΄뤇�n\���0<|E��#�6�*�S��A�t�ܦI��!=Ǎ��,/LqPnU�Tɴr�ġ��)5��R�4|Ĝ|r����I�;��A)I��JJۦ?l��ե��σ����N*�M1O�_��'�ajւ��	�
M�$֎z[��a��;�e�B��U��N��ؕ(��ov2����L�x�W�Yq��>/s�_�Vq�W7�f	��_���R��2C��7���i�	������'��'�Ē��+�37�TL�,09	�e�;fU�1��r7@��i��^�u�Ri����p{"rW�L��k�>�-yKw hmū;țW��9�ꍌ��c�����������/�oMW4� ��l[.���d<g����!k�7�7J�P��)�O�%�.[ޕ����Z;JK��b���0/���j��=���7ZM� r�y���g6A	;�w8�E!L��W��=����B��o(J��l�a�VK�"Dc0���yh�^��&��,�͇�6�:� �K�_e3#"5мk-�5�"��ڒ���l��q?�fN��f��
4�1�X�����S�k�@���Y��\9�N�/���e��3.��
�Q]�ӊ�2x�=	��>��h2<���q�	�')jz">�H������?�
L܂�e<g��氽"�"2t0o2��-�����t��Asƿ�a�-c� �껻�࿩��E���Ƨ��T������_�H|�J�W���PQ�&1�E*�#Y�b��%x1Ŧ��G*���S�*t��*B/�4�e�wt�44��)���Y��� ��^5�I։��I]�h.���A����~
l�X�R��H�0�,�,��)ڙK��3�kIgD�h��,SBB^<���S�W��\nCD&c蠟ωtB�-v�{�{�gr�e\`�znW%L����"��+&�~�1���
��#�CJnpbk ��g�����Y�0h!�`�ߔ���~�F3%\��"u� ��_��
��.�E���o�xM��B-RR1��%?�Vlk��g���_�W��zFt�oͥq�M�p�9�9��֊��+3�$��"o�uD�ڜ�UH�;��[.p.�`�.L}���Eqź�����y��1�->��R!�ړ:�����F������u1�?#�~J?V�	��2Eu�t�.�B�[��`a)��cMhc3Hވ�$���N�mZl�j������OP\Z�dm-�?྅9b�ﻜ�JH�C��/�3vw^��ʐ�8��Ǘ�r���p'G�>��7��:�T�q���ZA׆�\�t�ό�X�5�Ɂ�+K�[&VC�n���oI�1��������,�u�Dj� �!T����7!y�bɍ�x�/���}�� m8򋨷��%�w#0����ө�y7�W���� Y~�,��J�_���:�MD��pp���Ρ����6�B�#'�0�ʹ����Z�7>�P@t�A�0U=K�E�"A��MW���U�X#I@'�C��fJz���)�iN�����S��72�/��� ��ɱ!4g�*�굮��n�Q�U������x75�<q��Gܖ8`M9 �"]:3�6��	6�(�%X�m�f���|eD�0JMW���ō�+��q�}x�8��NЙ�c"�f���]��|_�GC�g��: �y�:�,_]�1�}�HYOGo�p���2��Zػ����Vgzt�@!a1���~ d�KQ�l���UY��x�xy�����{5j���.��m>g	=Bh;Ա<좾p8*LEr)�h�1X�X�@�_�Ƅ)��I��^9���I���YU]��Xل�9�K�
Z��� �O��\<Fa��L�r�ņ����w�n�Rg���7V������R�+Z��#p�/Qsyi��$�(��<R����eWטw��:��d�U8����h�>�]���Q��ö�0��<���Yˉ��Rs�|���TQl��]�X�?U�$c�+���z�
j������5Y�f�O�B\Jyw�-�k�<t�e��ڂ�b�\�u,^=�����p�m��0?	X����Gq�@}��~�o�9� �
|�Ѱ<hA@:ة�z���6x�6	z//h!�� ��a&Կ���џ8a�*;q,��< ���oe=|t>���Z	��O\�m�>4��̂��D'�ԊZ\[ð�_���Q��-�#�"	�y:d2*�.�
��C�&��_&�+�����tz9GnlجH{�����˧v�TIg��<y��y� j���P�Y_�8 �7��%W#��Bk@�?��(��L��Q���Bӄ?�(��֖2bez�>~?��\�<�W��=В(�OYw�L� �	K9�J<�<7���A�x� m�*$�
������L)<�m�]�ʆڗ�����=t�7�VZyx��#��Kk��%rTh��opi��%4%+f7�#��5ͬ�f��dK�C*S��d��i�Jk���Eܫ���@���&l����Rr�YX<m��r�������nZ�2��*�cuEЂU4��A�M[��.G_U�"����n֪�Rp�/�wU[�~ ���r���Ɯ���FI��6Es�K�V$	bi;����,����:	Zg�49��_"ި�wd��z��� _%�r�'u�9���n��=�Zʠ �6�j��=��Tܾ;<�=NR�)z�\8�W.��ͫbg��_�1�k�f<kC�]�5���w�EyY��Ǽ؋�Y1Y+���R��b�*�Ծ�	8��K�þ�4b���h+L0^��Z��Т���ja��ڊ1�k��jЖ�/�7qhN;"�jS/0�%�Ma�>�����ָE}ԧ�Yc/�9�VW��]O�J�0�O�Q-\WĊ�����Oж�!K�m͂
X;Pr�/�~L���34�˜��zPʞ���+���~p��7��Ȑe�n�E(m�|�������<��#%c�?�Z��ɕjc��`�B$ߠ�������}��o���
���� ~o�߱Ӥ� *H3�U���ur��G`$Wj��X�Go|0�ek��(np�:���9�:���'|3�ޕ�+�2;Kj��D� ���$��]_����r�}��Ȩ2B����mO���c?4-oU֘�BR7��.~�b:J�{n��49Yr�cۑ��ձؗ���X������f`�����E��{��!�%�����Ki�| �kڣd�~��;������RU6��ڳ�����u����������p�BKw_��M
���^�bo5՘�&���JN�E��m�ȃ^�C��֗Ǉ�d��}���YT`���*��zR���J:5u��b/-1]+K������4A/#�r����v�ѲX<�~���zl"��+��$���}����m�2��J��\��kTﴬ;4���čC0�/̗�b�Q�-��RGN����� �'`��ƚ�X��A��s?��8��":����ȗ�;�V�33�֞�.�ՠ5�>�k{*�*c�Vo���<�֐�u�|��wm�l�1�FzY]�~�u7�d�]���>���]�~z�gpԠ�u��K�]� ����KP�FD�3P��,p.$�`���ʶ�X� �ͽ��D�ښL���wy��*�U�d
��� ���:+�g�T#�V�V�� ��S�*F�=���c�C��5��c��(�[��L� u�n/��W�����k���e� Q��P�� �~��{���W\����-aJ��@��-�%|�Y�(�ٖo��q+�n<�@	6A�Ϥ)]��L�d�pb��S��������FN��_�=vuA�E�7n+���#����0Q&��͂A����0~L�/�(��uo�?}��hpL��)�x�0�f��}�J���D"� 70�;�l���K]��W�x��n3z]Q��@� mU���eL9�I{��c�:aۉ��ݿ��N��7o�N��l�X ����E*��$��5�B+C�o�{�Z??D�W�E>r�=[�N�w�b{}a΀H� v�.T	o����L ԯ�#_K>G���~�Y�h���K�@,�ai��_Ĕ֖���tD�6��?��C�N����
\w�ϊ�r�Y��4��k�0!�#v��$�
�~��Ic�"�9���UP�b���u� ����=��+������&�j�Id�R��=&*p�_Hm.�0%��Z�kY\:|�ΐ�jn��a�%;��f���8|�'�"����JP�c��w��W�C}?��[麱�mM���~�[-ה9�Ѭ׍��_LØ�ۣ�$����'����9�q ��q�#�
�M�g^[VV��Δ���B���Ĺ�~2��Nm�T׳�Q>c�����Oz�	�y���S����\bKc��&w��Ed�xCG��7�����;�?;@��2Xa��Q�ˁ���Ñ8�1V-�#�男 ��߉5.�p���g,��(��"����@�¨��w�.5�جֽO�˶"�y��)d1о�hh{X�q􀙩��z��q�NWQ�]���7�^�Bޙ���*�UŀP\��o��>v֟܉ ��1��K��ᘟ	w�)�:�(��_���+ms�,���O[��������Kh	�M$4]1�<R�奮�̅�Ak��Je��{�]��3��+���'O�f�k�D~�\��lK��!������d����l\�� �4yƉ��3Y���o��q�_9Z	��к��o��i���Yɒ��p�7�C#�Ti�S�����~}�*TK�}������b�~7d3�[��6t�R^�5Ӟ� �����=��$�ܹ���_G�t(��cXX[io�a�����z��F��k ��b?��T��FJ��]
���w��Q��T�@��(Xqb�� �C�	5 \,c�.#ig9T܇��C,Uk��6�+NЦ���%���D���N.����cr��TQ�e�ͻ��b�a�t����8 �ƫ~��t��H��ZjN-�\���۪���I�h�q����oה� y��	�-��oMa�ia2zORc;z����9�%���D�e2.�^�2 �3�� �p�3<%Y.�)�-��J^�T�ܫ*??K�QO���%|wU�u�u�}��b����.���&e��Z�J/�i�����Y�z�h�E+��yl�B0z��{i��-����pz��1}�������� _�ʃm��&�~�g�1��-VET1��Eb���K�C᭯�E�7�X��ٶ�R���&"����������إ׻��Y��	f�k���
G���� R�num����:�89�� ����ձ�4L,ʌ��0m�������9{�)O�{x[�MA��sQ$�.h���N�x(�+�e#Sm����	,��R��:�<�t�&�3�zǁzC��xD�;��G�<Mfo�Ĕ��k������*RV��#��� e�5��B׉ef�̄9�Y1QR]�%G�5&N��[|V�w�]����|I���~�[ӆ�t��i�4���[��HJ*-疌�������t���9�1JR�4�q	�(G�O��{
1W�)bW���!�C쾝�2Iv�Ju6ر	k4;�y�!�HiO!g��M��� ��rb��j��>��ΚY��h:*�,�L	�*��C��p�p��^q�����A��#"�q�� �t�yIg�z-QA\	��N���r&����+q��i+w�^ͅ6	��e����y}QtD�nM�Y+��I���=�cq[2ꨟ�a0�"��P����5�|6+��?��8��e���4���p�}��н�E�;��q�^��o��h�����C�#�7�^����R��z��Ye[�N�ѡY�5���p����
����E��3/��
bi5n&z0����:��$�bɉO�OƯ&W��:i`.��rᇮ��B�h����Ɣ����Gs�PT�v� �r�p�[���alg����5����k�!����Y�	��H�;��Y�"8'��|� �e<Wy	�ٕԼ��lg�h���N {^"��5�6���K�� �k=!��8H��,Ŧ[��AU����R<:�n�@�\� �I���F�ܡ���>4��{B���Á;2F�u+F�k�S�P���� SN�^�xV�r�̖#���@X�ej%��j�e�,,�T6���J)ZrK�/��t��E40	ھ:��7lA��:����A�V�n�!Vc��%e�ԸN8ɸ�r�r�>����0��c��hT���Ja�G���"/�m��`��pnv�t�+��iF�� G_0�Ʌq�_��S�-H����GӍ2C�w�Z�C���I�:1���i|��
Wr���5C3�r*��>��N�S�<�Վ�A6ZI����YވH�7�ɐ��"=܊��S��iÞU�c��*f���s#�C��(�>S6W��2���NX�_F%�1Ws��Ҕ�p�nu0˾���o�#���g�����1HNN1�C28:@;8�\�&�Ӫ�}�eM��F�i��)z���}>:�)�p�_�Y�����]�j��/���x�Hu��۷\���7��6��ә��� ì8�=�������?l|T�ryv�B����Z��z0��w�}m�x�x}����=��H��0O��݈w�|���ϩU7~�������*�k�b�N�D�&����ѐWY�B�ã����i8'�M�{zS(�R���;�Ѭ3��yf@�l�e��QXe��
�qf:b���\�+��o�T?M��Z3$��y�hr>e��h�N~�Uًv���Z�/�`�)%4|����}\�� ��&0kN��Q��}MN�d��#N\ߖ���LN4CPWD�'�j K��F0�[�#�p��n�Ի����.�`��I��Y��6],H9_��^�#��������e���[���7��E#M�vY���č� �o�-�V>�cR`�	n�j���mΘ�C�3kf��]v�g3�LB�����2y��TZ2^\5�_���`��$���9���Z�b{E�FB�f�hDn`4R�{���u�xX��b��,���%�i���:�V�����A�ú��#���N����b�K�0�l��ԂW�-X�8|Q97@�`��X,�R��_Gy��}�%0؁Q����\���k;��@M��"ݮ�/�N�q�?w"��t�c��4qw��.d:ŕ��N�:d��t>e�*�p��,p�*?0��NuAW6Y>c��`T�������j��Yudw����9��`�_��y�6��j����Aq�f�����n�z���U �Z�6�h%�� �/f2�ǲ=״�^ۢ��������H��T�6�n�"�b����Q,oDi�z*e�# ����g�I��:9��̌SP$��j�?.�>��}K.|�Abk\t���0��{.��T���s�wU{,�`�HBf��|^��O������2E�m2Y���Eo�l����&ѫ�f&8g,:)JJ��+��Ў`5��;s�b�� ��*�bQ�{c�H=߂O]�p^�l��b��VGAc\��қ���eKݥ,���{���Ԇ%e�&��&�<e�dPQ�+�iN��8�"��Es���cvs�ϓ'0�i����r��Q����wZY��tB]'��!����`�0q�)UO����0������F"��(VD6�ZX�Y�7�W��7�(����U�	�M��%T�%lE���춟#DV�_��z������Vr�VI��k@U��߳.c����f�L���?P�����3�,
����S�:�yU�	���)�ŷ��D�`�.����Y�V�3Ҡ8�����1/�t�W�H�
"�\X��gAw����Q��+��7W��@����=w8z�P�]uGT�����������l��bv`��.��}�_bN���A��{�@y�r�����)VR�"��&�4O����_u2+R�D��$��u�����ʹY��&+��ꄋ}%٧1@�'��}#�B#;C'��Faa�Z8����R\_��,p�����MV�ݼ�1kc�S���
|XLC0����0@Ar��&we�/3�r�lm�>�Z�7�UW8��T�}j����r����u���lD��H��jR�����Go�&D۞vDn�BW<��y���v߆c�å�:�Wa����t׶��j�4���h��yTb���;�<����}��G��i/��J��_����D���t�b��rY���r���f&�	�Ao���(��K�d�3�DF.�_��M��l�����Z�K��v���.a$�WN��� ��F=��2I	�U���P&1��w�g��&Q�����l+��P�˛(��TS����?	�֔�H���Z���`�$�O?�L9G�k�-0↉s_i�"[N꒑��<���9:����jZ�ޝi9���.�Mce�<A�
��<_h�c�b�1�ndɲ���8核������L�-�T�#���6Q!H9����DK�	�j����K��{���۽��ݑ��L�[���LuU���[z}���8S��K�&fn%��i��vmVU����Q��h�;�Ն|9���>����?`y$ڝӖ Nkgx*xҧBf4��e���HN���N�"��+���ŷ� ����#�]�QV��{�,ܨzz�M���TY(��z�c� M��F�+��Q��'�<0%�`���tH���9/%�[���j1Yw}Һ1.��I����E�)3�~��ƺ��1<�H&�����R��'�U�Z͋�]�S�{�&����� ��^�6Bk�n(�h���V��GH8ݭ�y@F`[zv���H%!�^�TP�'��w䏾��7� E�]5M4z��0��=1����)�JFF`2ДK���{54�o����>0�p�`3���Զ��/)�o���Ŭ�����"g�+�a����0��¼���+HG�x��Å_��Q��g�g)��eI�$.�PJ�V��
�MJas��t/��.�a}�jߦ���ʦREz�E�q��Zv���6v���&
�V>H�!��T�JR�*6qur)�I��c��ƀ���AA�z�}��&�T{j Y���~9�raL=�]W����E�(ha��ROd�}Fp#˹���b�w�f�+ ei���n��UI�i|����3B|Ck���F����h��� �J�ɀVuW-
���aD��!�d��ث/I���P�eZU��e|\q>�ʇ��"��4����	�t̻C�ɀMi|y0k���_r�-bΫK��8���k(�����yh0�iq�BB�w���p[Q�͚��k�y�A���m<T�Ed2�g��4�hٖ-�ԣs 0���w��QA4�L�o!�쿴Y�&�(8����X��"a�3%� ��W�z�����g�]"dt��N�6	2����C���op̮�jm��5\�L��C�L��ujL���[)�����^�<5�/tU�V�3}0�	�aK$ �7ȫ:�*��� ��0�3��T0M��2U,�b��Q�RCN������a�H�������N(���[B9���x94�Ka5� g��k[�
L��3�%���2�[0엶.O%D(ʹ-�ڽ�U�F-�H�vFƃ�^��Fd(@m}E�����S����)wD�f#j
ьWH�2
¼
�H���I�.�K�ð1�B�,�ԧ��KU	��%�e����r�)�Jm���z[�?��3�ɥ�4�����k)>�x� ���2���8|�S�5ZN%�!C������>�V���f��w@qFT(9f�	?T��ͮW`3N!��b�ۥO�+�Ax}ү2��ȓ�4��9"��ڂv��T=C��N8c/W#J|�6��o��J�ɑ��k�p� :*s�����?4��*�vc
��������тa0}���U^��Ϝ�ˣ��ە�X4�lԛ�Ľ�Rmn8<��J�&-�e�\,��F�1C
�4�vד����X9N��)�0�����cAG*���:��-���W �bu�G5���%���+Q~N�w%��tWH^챼���e�MF��9�^Bs���޾9y�%R_CW���+
�7�����h���v��bz7�Y,OU�SkXӣH�\�9��}��G��U	u���1��\�������j�(P��d�<m�\ʒ�t�q8(�d�"�A�#n���/4�V�0G����#$	�}�E�94�qgH�,U�FZ�x%	b�RDUM�.�g|q¼_aGF�C>�L�hd���C����"�S�y�ό �#�b�lܨpy�{�||ab	��fI�H���%E'݌���@�vL54a���|�Ǳ�ݧ�Dt�ڋ�IdƎ�f_�H4������wZr����4Vm���Ab��coح��?i�hPqf[��'+h�fY��1u B���J&�-�ȐfEʊ>���o�o�3�Tʳ7P���""@�'��M�"-�^��#�
��(w�C�a��A�"��b-d���"�"�X�3�
$�����?�A���aɮ�Q��IR��ik��1�I�	�Y%�9+n�~���� ��^f�.�q.������ǫ����b&�MЃ��!|�D��{e���i����̬��~�,�f�'To>z1��ZU� �*���Z��g�n�)�]!l�_�۠��{�<h��н��^�9�äJ���z�W]-o�eY�i���&1Q��Y���g_�B�m�0������c�����nѳ��B��G�n�$�����c�ԑm`��Q1�,@�zb�?p"^T�iD�LHr����&9:1e0ʼ�M'OF ������$�����R��({4��t?"�'�F�Z�)���R{��9|�e"-��o>�ѐ�(��X�n�n�jb���'"������� ��q�8�ڎъl��	,m��v� 7��>V���R�󑖇TE��.�r�C�,�8���8��9��A
��#x�>�W�����,{+��ݬ��o���Cא4�n�SQ1P������9,���hKk^"�^ÿ��Vΰ�d���*��?�����V��4b\��3�1�@�*�AR#��U}�F疶`H+��$3! ��5L��MtHX�d������I��JF
*E�+����?z�+wY-p=����AT{%�I�T�y~<�f�\GY� ��k��� =on)=�$۵}(,E�@�b�W@B�/[c���Z����ZP��>1��d�TQ�p�oA���,�Q&M�\��tX"��RN���U#��Cw�_ɲ��ߊƃb,�=H��|�g0(�[][DI�j��Z�,�`8�����^1j�Vz�A
(�G�j�ZD,�S�S������rz?[�3"����A����-Bpv��ubr�
~jyS4:VH�	h��e�t��yf>�s�CXk���!j�yи�aA��L�>��Kv_y��;�.7����k�w=�PjEJ��a���%ѻo:��(BH�%�����de鞭�4���G�1i���	��m�ЮP�����K�\����$�Q�<Tq���j�6{�� ��񙿝��������'��ߗ�����FZ�R����\�V4��R�~$�C���5�MFOvG>N8�� �#7ɸ��c�����x��A���,:t��Da�i,$�;�Wt{���G�lrȬ�$m ܘ�����3tŢ���U�^�$+��໯�!��GE.���Hd�u���^��y�1�}}h Q6!�39S���Z��^��`|V��&{ ����UH	7�1d �9a~���y}~�{�ң��|��k̈�O.�W, D�Ço�Gک��XJF�/N�d�#+uE��p�T�=$�oOw�lț� �T�+$s���\Q�Y�e�$|~��Y���A�Bw�c�"�*aZ5�w���K&h4���c��:�<��0Ff)���µP�����lJ9_؅�3���(X�I��$P9����D���<�̎������\v��-�6_J84�g�3x�J� �a��J����kE�4"x|Ϩ"��I���|���՗��cb�^2�
��\�a�v���@�C�x�ج';�~�����/W\k��	��Ô�+���;��=q	_V[\� >�^<�)8����ܓ8�q�}�Ú���<����8��L��_�q�J���1EǸ��ap�'h�wGe�M�d�!~]��f�^���_���I�tv���4vc�N���f0��1�����R�
�:o�2@'�c֯y�5���h��T��i0�zS�s�4�E|?��'�U�"c.kQ=��v���[b{�ip^�[j�?�R1�]p�Gg�1v|Dˡ��;���-_~��>�0��+���$��94�Dx��m��O=�ȓC�ZK�])��p�1��5�+���Ū��>�z�B�F/�$��2���n�Y5Ɖ�4;���e�h@pn��tE�4`��8�aY��z��ʭJq�m��� �o�Чn1,,�|�����Ie�+q!��]���Ɍ5"_�_�mE�ew�d]o�S^������7!�*��n��HU�$5�pRiw��_�ͽ��VK�x��X*ɣ��K���Y�����{w�| P�������� ���K�;�a	s�$�&w�X��(�$�I�=�"D�ڗ�vS9լR���bK�?b&[r�tCTl�>�#�����Ι�F���>HtCw����3ks�y�#���;Y�?�K]z�c���U]����U�ā~��kj���!u]-s��f�K�8���t:_��w6f;�4�/�@sH����%��.���/ �n�����(y ��T�2�~�T�����C�rf��B*�Zǃ���S�j���7�u�3���2\�`�����xx�Y_��Zo%����(FH��0�������k�������VM��y�nfc�.��Bs'��x��5gϰM;>�9��j�묙_�6��k�.EF_o�:A�o#;O)Mѫ�!Hn�-�R�"�2�+H|�t-89�t��M�g�o���<k����p)���8�E��FOC�+��˰�~!
��7 لj��L<ZM1MŔ�ro�'�w���'���Ӱ��� �;J�pVj�x���?C���J[I�ڵ���G����^�J�f9b�F-5�
�:ǒ�oY����G�3�/�>�����C�}ѵ+~��@܌'&ﶈn��O�g�fF7y�YVt���,�0�br�-���r�q�}tT��ڛ��Q��P�k������r��'�T�zq$��jÌ�i؃��6j�m�:�T:3u<��N+q�G@`Ʈ!��U�4%KN��"Uq�7|^�U����%���{j������=	� �|�b�G�����y�cG� �=~e��	��7;�Qd3��;ɛ�N��dĵ��˻Aб��8�Km5��
U��ୌn�t4닎|/��ݬ�<��M�n�i�6���\���s���QukW��W��%��T�}ޘ�dz�&l�Ջ���:*;-�?�	`�w���l&fZf��}�)����oQ���7ʩR���bk}V��i"�D���ڲ~\;~����_4���;z���Ɔ}����M86_P]b�O���������9����BP��*��^�X�(��x����� ���'�E�<w�����c�	���0Wz�@]·����x��i=�@��7��N?�9�wsn��\o`r�R���$���%�����vL�h�*�<���<�f�m��P�S�C�
��NR���
g.�_��+�	��Z��%F��Qݘ����ʃ��>�X~kЮ!i���tR���7Y4�E}L����Pc�S�M&C<7�#x�̎�]�
>��Veъ��̽;����[�'�?C��f�(�+м��b�7�w	k�.V 5 4�%�{k��֗P[�&}Mo��;u���(��mU���#s$�j������}�^��H�W�f����WƁI{��U��Oz>��;$U���K�3HlAc,fRB�k�q��nd��i���tИ�J'\�7��%%��^�\������N�s��^��iU�2)�
n�)n;2ɩ;l�	��(x��'}�A��,��/��+X�a�l� A������t�xHG��㳇�����ު9�ς��K�sj�ScCVօ��H�3 =���W���V.�^����Fz�g�Ճ�:�����/=�4Nȍ?�g���B�<��fR�"���LR�?����h��gn4���}���ĵ��d4H&T/��C�8�N�r��6(}'T�O3�0��l���ڻyfǌ&0d���sg��*�\����]j!��*@)J���4G�P/�5�� ��N~؅&�:�P}n�0{���5��Y���k��1��I�;�<�����j�� p�����)E$����o�͊ �#!���)�9VY����,k�p������֗z��A����ׄeV�@��m7ѝ�:j�?4^cr��?t��;�5w��u�'�%_�&���3����q�:U|�h0`.K��L��1Y㕃�kZ���yK��(s���C����z�/D��u�¹ט�+�]�(jS��u�kⶲ���I�p��|N`��r��*?۲�t>�w&�6:��`A��	���"j���cϖ���[�¨=�����q|љ��M�����d�dL�B!t�}x�
�r�׵���V�ﱚ�ۉ��y�]^�KR5j��g��z 
h~$�Y�2�a*-R��n#�jK�fz�v�g��m�� ��r�#M��^L24u����ɧG�g�_z���%�d_r�� /��<���z���Ç#�틽����Uqk�N G��^B>R��$�h��L����q�m$�m�����j�]����xA��0!Y���}�:z�\aE�G�X�����KD�����[Wr���9-dw:����li����^u�M�ᔚ�z`1-�E���5�
}���ץg��r�y"��:��3��Lo(��M:\6��v�uD��<����?n]���rg�0�N����]������_=X%�����>�n�e�`@��_��qP�\6ӣ�(�
�2�c{;*� �r� ẙ������6�Z�>kꠘ=#d�(�M\��,�ݢ۴�K�G�&#}nV�R�n�M��Ba�}2�.���5-=ÎtF0��Mz����Nuu�7�6���Uv:hf��'��ixN����Gnj��2Ea=�?����Zޮ�?��A��T���+&SƁmE��R
�5��Z+�}4���k"����q�]��J��cg����~B�4��zO��N��:%>+	�\f��ͽ�3E�l�x;Ʊ(k�4)'}�S���
�֯c0|�����;�ag��{��@�sL�_zc���B���*�v{f�n���
�'C�E����XR՞O
�bk2�.1��cQ`ݏU$�YOͲ�K;5,ō��m��VT$GT�ų��S?��k�/��W����ق͢�j�H���֞#�6��Ӭ2�J��u�fӱ���Ͳ�AJ������ؼ@1�뼾��)\C���l��><���ƣz�5����40��N��j~X/R�Ƶ����LM������uԮ2Y#뛑B?�7�m���VV6fR�����O
�u�21R�v��В��(=|�t,�0X��}��|�?횣��L����4klQ�"K����dk�2��ϵW0��\\�*����/� O��W������F�90�5�bO��ߚp�Pl�G����ҍ�,�mn�wq��)K�]A�K��VGs���f��o<d[�-�G�ʤH	D���^թ�r_4]CnŅ�9��/��������a^� �ꇥo^yx��(�`5`��W1u��>
9��G�<d2��=C��ݲ�A�t2���/gj��v�
������iبxT�c-�~��;�%����*�����Q��U�N1NsB�h'�2�� �9�`��Ɍs�W
���l��/=�`�	4!V-0��6��Y��`�c�p/[H*\�]aw��]�
�S���4�g{C�
C��Y�E�)lqe�&�N���=�|�jE$!ɓah���1�w��0Jd��T��BX�,���p�*���5b���&Q�^��+�%�i�����ifk��
v$�S{l��nt�4q�GK⧗�C#�
�[O�qj\��	R�?�7�s잏�3���H/�)�V̓h��GD�B�(�kT��q7��)'��,!��[����r�D˪�F��ҹ?���P��;�ΔL��ޜ=p}u�	���P�S~K;a/����_�W���O(0�6�Ձ��y鱈�Ff�x��Y�_(�ɐKd+ۙP���K�K� ������BO��yѰ-"kwZ��~�I��G�>�q�G���$
NH�`�.y�ɀ3�J]FZV��0^�L���YP�,��Y��5�G��$T�C��ǋ���6�$_�^��3������B[��Οoe!:j�7���6�E9D\�(�_W��I�L�����G��!5wS�?J�\��m�c�S���/3Pqi��������Z������*=C��ODu��J��c�v)!�#]*�ޮ�y�a_��Pm9>����i(�·��u��z�(:,r=��Ē��
6��v�k5=9�S$�Ŷ�-�1]��@-�Wj��Ѧ%�5DJw�Ma�b}���g*�kf�Pr�ҷ����X�@�&�m�k�A�DDv8��eXJ����A��w�}p���a�yyb�/�}��G��LY}�dL�j^�W�^���IEA�ob�8D�37A�k!�~9���Kݗ�UD��W�j4�0<���@��n�4�-�0r�7\���i�b;��Q��/?�M#dh���}����R.?հ���*�
Sǥ	O���[��Ul�p�>A��HLmq�]]����J*]U0�,�g��[@���do�P3A�]�~������ޒ�㣝n(�;P�&��X+a�kW��*��,���͙�������c�v̇���m�}��^ȗͶ�c��=~�z�)��J:�40���Jռ�{�5|�Mf��M�i�?F�(���}�����@�ӹQ�i�'_��fu��{���Q�x��^`'���ص�u�k��gl/�~,�N��hR)�˩Nt���>U��uz}�k���]c�������{��M}����6��=��"��X�B��`k&&�!o ��I�iG��
��[
fT��N�`�?�+�"���<	]����!^�ef��Z�߇��L�ŦJ�:D�F6D��s��0
�_�ssY>k��yX����3ޙ�o\62�s?M�öy�]��`�@��яI�?�3��� ����y�g����l�]4FG׽�$r��o�O�9�"8�n�D8d���EP�����3�����wJ�lsA���&MG1�LʃY~�l���^�t��V�#*e����8cqzP9�W0/��k#�-v�+j��[���s0[~����8*� ��"����_�'}�PI�����1o��;��(Vz�N���L��?J�Z��d񻷨�=F�����QZ�D B�Xb�����to3�n�;9"�Fo�%�YP�m� �!�g�4k�w?[Nt��h�����[3$e���~��w"u��]G�qs����K�a�����l�8�^�@�Z���>�W�X(�آ�%�:7@J_
�{I���u_�2����~^���>�����>���>�/b!���e͑4_�9n������r��տD0��$��!d�W��oAՌ�S��Ŋ@�t�%Z�e�k}aϤ&��<��#
i�[+F�ZȇB0��R�b7�C�]��'p#c��# 1��c�{2�X��(�������\�������ڳ��F��dؙ2���4����_E� �R�ۆ�\�%�ĀZ,*�p%���Qsr�N��O�e*�Yո�E�<{��z�D�bkn� ��_�������%��j�� e��3M^&;�%��%�o�sC��wI,|�u���_&:�:W��Z1պ
U)�n��LPc�
S�:h�~t�s ��"�"�H̼{�]]8C����ܯ�
o�!��YR���*v�#]����(u�ðA̺a{�Yh�X	���=O0xc\�/Sn��S&�I(o�*pk�HR��/�1�a�F�*��ǅR��#�2��-	$3;��l�`\r�|������TT�u.�ּ:QcT�y�ЦY�<��I��Ǎ�d~�;���~>��S�����w�+�Y�k:�b���/g8}G�������!L�<
�#h���䛦�ݯ3m�)�"����"�֦QQ�C���]�M�eH��M��K�ϻ��C��4��!~u���˿䑘�bhdx~J��~�&�m�g5�6)�ǒ�� wP���@�I�������!�y�)�[Oo��#���v����bAJrL�+��,!�B>K���X��db��R�����&����I��kA�-ol�!�����S!8g�C���j�+)�+��5Re���&<j!���sS *��6�7?��Ge^��ۻ�w*L�u���H���
gȲ@	�FA\����ʷ�d�>���6��{l�x)���p�
�����.�$�^�Y0����ª�����f�8Մ��V>�ƹ�A:�[�F<���4Q���2�X����8OIU��Mm燛a2\��&=o�Y&�a��1�Me��R<W7W�`~��7�"�/ܲ=������|�*�I�P�F���ջy���/4�,�ϳ�&�(-��l7��޾�WVO�?�]��irJ��9���_�$mׇ
;S�m�A�ŀqD��t�[A��Yc��F`$�E$@��'�W�A"�ܺzB@��Ÿ���9�PN�i�̞�z���{�(ڬ�C~��-�\����wވ����L����#�a�;$�JȻ@��U�ٜP�/9��F����i��DR����s�r���r����ŷ::����� p�e;)7C�ⶍ��_���o�3X�S�ɵ���� �7�s��=Bf �c����F4U�c�2�Y�@�*zHR���C���B;g(����lМ2]��9̫����������SH��TƈΞFLX.��Mfv��t�zPX�;WrW�#��+�N̕�N~DV��?-�^#�F�Vz~=����s�@�P
�/R��k�-�(�1����V5?9�F��ךs�"��W�յ���~��p��<��(�c���F!1W�ח��1A7j�Z����_5���7���S(�� q��+�o�O�L�i�?�����%�%Sb6/Q���W�vnT�5����$gtiKDPR>�s��u������*�!�b�y��9Z >=bN׺c;\���w{þ1$�q�XŝmW��Ͱ��`�ɷD�Ɍ	��I#6%�o�9�bי��U�3�
k�M����e�\�D���X]P�N������o��Sb�˲2�
�+���Sj�J3�h^��_Y��_���h��"��&y�G�ɺӎ�>���.F���u��B��^?��ԇ���L6c��a��,������������a�:�"�8�F�s�=鉌�&�$���#��ݹ��t7�g|�`YL����Ճ��!�?W��8<ɦ�/����F�v۲5Ez�.Q�v�A������=ץ���4�ť���v M�6JC�+�����,�8���p
s6|r>�"�Ix�b�ߍ`�OO͜����s/�}�.����λ B��deL�o�W�I.��^�e�:�����P&s�e�T��RB�5n
�
��I����.���g:�l����7j�!=�l�9�q���Q�g�����qc.O��?:��s+�Z��O*X�(`vĄ	�n4�h��׬��R>�I���csm��턾�蚚����6S���-+)��%�i�u~�$��_���qǴ���uB��̤�����U�����m�qm-"��!8�)�(Ñg���8�r�Y���p�A �d�o�>�!��/�:�w�ҹ�y;tA?�q�M�#"{�8���!�az�r�N��h09��7�Jw���#7�L�"�hlPn)#˫|�vh��U��ŷ�@��9�#Twv�K���8���c�5���A��V�� Y��s�]A��!�rl����%0
�?@�VZ�7<�-������(��<�Z�Ͻ�=�t��4��&�O����"�\ETǫm�����C`Y	4�0��>]�i*��w�BYQ�:6��y�/�5n����U�E�e�\3�y(��C�!�۷�ݒB�5D8��2��\���Z(���<3%J�D6��ܢo��iH�(~`�{��GfU��%� ['��_��^3��[���V|K{�%�>��;��zOi�|����q҃eE&�����SU�}�֐��ed�ƘPXa��<��?u�����Q���N�Z���i��.�L��x��NW��P]��xp�.��!���D�E����;M��/�/�Gu]�z�w���[>�O�Ϣ��n�r1o�OI�o��f�{l��� ����峄�
Sڊ�d��g�\��j��x��?��Hߜ�B�~� ����O�	>�ŭ��6���)ض��miWL����Q�[8��L���;4������88�ۓH�����Z��p9��Ķ����o�s��ï`������0t{��K���/��|����3y������ݗU��� �G�j�O�3�cˎ�`0�j�b�/\��^C@�
�D�1�]�b���XTg��v���Ncp��:�i����O	h���F���3D��V�zT4��)�ٶ~��5a�$� �7�t;���
U2��m�2E`Q�k �[��8����r`��oCqt*�p.r�H��1�;I�^l�kz5ȩA%PO�Eȧ��	����N����`���HSlh��:}�@��[UW}܆�a+��OP�h�����}�E�jKⰇX*\ë�)��q���+x�	��y�<?Q��%���9k9����8�W{Y	�#]�J��.m��A���.w���P ��p�Oe����5깎o3t}:3G�W1?�V�V����kPY��*��*hV��x>P*LU�V��{K�۽M@�_/�+t�1[����,_U(r��#�F�RC��5�����I:��"�M��Gϡ��^�\�����ﷻ݆w���u����j�!�;���w����2Q�I����yA0�
ms���m�0뚉��]�os5�S���p�P3��z���emHIc>�dV��	�L5������J�!$�'N��A����a�^7�VFe��UQ(��]EִYnK�4���?w�qr�v~;|j��)�n�`�̈́��&g��`~7zJ�1&~�.��t�{enb���n�1H�ʝ��UR��qaF�<�nM������z�H��	�v��}_k�������7"��jT<��`��k������6R�l\��pVY�m�(�Cw�lSb��L)����_=4?�|����,Z�C*u��>���9�#�,i�Z%^@����l��mj���T?�/�l�LP
�W�wӏ��O,��F���`�j�j��x�ٰ��(��K#���T�P@E~+�F�Du&�����
��N�Un�n���E^���v��/��3c�6muŜ�D�* �du�)j�EAeO��ٮ�t�kʓ�ۄk�>������R�Ϡ,u��L�Yq��dUn�d���H�e�q���ۖW1/곞; Ɋ[QH`7� l��>���O.rU���s�����[���H�3�w;2���
��nE�� w�����Y�05Ec�@�a��g�T��-tXE{�(O]�6�Hݾ\}P@�&�R}E�,�Dx��Q�������������WwN2�qfS���6 sXJ��q�j�l�98��Nfx%!7R�Jc��Z)p�Pv9��aY찐7�� _��}Kۻ�S��t�� ����2c`A�B�j�A�������u*�I�ݗ���G�"�F�F@0��k?�D�m�8(4eU��p����N��N9�P"�0��6�w R�q����hNK�����3Bx���ǚSJQ � ��kZir;L��r��a�%HEpj8�z-��ZR���������_Փf�Q���8*`p]��<X7����5�B��	��e���'�'D���S�Zf��r�]�rޢ����I0�yh'ȸʹ�r���H�Ƽl�0fu��`@:�RBO�e%��B4��H����=��R|-�����FL����P�J�:�T��r��h����+Kч����Ƀe��a�J0j���u<�G��yFB�#�� �$�S��c���_H
7�_+��Mf&t���u��,&.���I�w��NoS[j
��l�\�R���ߑUl�__���C�+t������t���X�ZR�$qЋ��T2#b��&A��O�/5�M�d�v���-@�H|��0����D�[_M�"*���S��_H���<9E�5N�,��u�� ^�bǚsr�j*R�S�ܫ�S0�ScĲ��;�DZ����0��O�ᱤ�4T�$����<ΆD�Gpӎ�eXX0k��zj-�&A�ieㆿ=ھ�n
˜�x�p��s&�BT�X�$ց��N���%O��ΜvN��A�v|U�M���}u��h�o�,x%)j�w\q�͘3����N:3��la,'5)I?�8;e�4񢫖y s$��	oQE��fV5���d��#�SV葈�0�h_b����A~��e�*H�w��	���#�GM���;b|E�4b��.���ٟ*��r<�+�ub��}��ډ�M�}C��`���=Ƀ.�7x���IW׈QK��sh�5��͆��R(�ֱ�uw(�9m�|'B8Gtz��U��#B@NA����7 ˑ����?є�������ܘ�T�x�����1��Ar�P����R$�)�|8A��T"��h�#���-�|��LpU��x�X�zZ�e�DY�v�K����S=�E����m����U�v]]�j�gW�>�I2n�I%O6B�Kܪ�#Ɂ2�;Jr�
=�!�&m!2`��J��7��qW�@�{LBf��,�D�8�*U��<l�r��������d��������ȩ]� 6���������� fP`�;���x���'��e��K<�5�ց ���?sL\��y�8E�C�ĩ�s���tZ,K�9Hms��}T�ݛe� �<�QT^�m,����I��&c��"�s*wE���[�ַ�D��J�����C!��¢�o���M��t��?~Mg�7~b����sP�W���	���6/�n�#�Gfj���t�x�J��DV��)"kcfCn��*��X�}9�#K_inok�,>�F�օ�ŧ{��g\�1�T��z�a���;sP���t �#��x�C�q�T�yi%,h��Ґ����Ʈ�a
��ڹ#F`��������� ���lCu��b��/�*�oG�P����fZpl�Y߶�P��Ʊ{�K/�u�
�Ø�s��1_�>��M+��Љ2����ɻ	�%�u�|��&�z�l�W�6[/��0�0��ٽ���W|�T�����`@O	m>b�t��f����8	 c�£e����M���x�1'=L��4v���9x�J��V��r.PA�6Y�<�0�gA�>���DK���u���W�!����\�m�L�\����Ku��~���
���7���p?� ��`Ճ(0L�Ľ���W��`�7T�ނc�����	���������Vĩ�$aK��h�xu���k�x%����Jɱ,ݠ���X��d�FL3��$}޳��k��m����h#}��!eA���(�\���-,��/j_^y�����[��`�ߕl8� ����d�~����	�n���^�AL'�Ss`Ɯ�K�����
6~�Ca��gU}�����5���j������Hdewe�h>�Js�>;zQ�fLw��o07YY7S�u!n�� "f@�t'���+����s���`z(8��-�/����� ��I�]�� PY ���)�@�
"��ޘ�=�1'�o�v�W���:��L0g�f�H��=��?�M��
�(�]�b�N��+�����%���%��4Ԉj�I��4G
�t����p��:1����'veҕ5���>�VI��[���\��(��C�p\�i��5U�R:ևw7��9��q
U�P,֫��&_����xW@cqw�b�~�}��>���3qز&}�,���<&�Nnx�um���9@@h��_e��kk~�Θn����Q�[�ę��OR��^%�v�b5:ZhR
a��֧m&7��o���:0��?��!OZ��3�V�1�F=��;Y>0�Y۴�(`l���Ykl������	<nUj��a���1;�0���s�
̮t�}R��1���AW�q�ׅ�˷I,�H�-�Ⱥ���_�J>|V���9@�a\޹�����n�r���|K�E
�����1�h�Fg���"�-�	1nF&�5�O1��{�p��ZZ�L�M#�5������Ax��@�b�W���	����٘SR,*���
��yę4{�#<ay"�b�MP���t�#�s��Dّ�6ؓ9"�em�dÃ�u�ߤ����P�Hn%�=.��$�6�N�x�M�J�|�KB�w(�nz ʨ�h�`���Ubf� �����Z�7Si��~���O�_�Ә_ ��2KtL
�~T�F��Ӊ�k���Ca���tp��Pޖ�u��/-���F^8a�o�'';KQ�I�\�����S��j�8/�k<w�q�a��W�pwҷ�˪�Z)�P��9����� P��F���!�	�z��D�w��j�F���$��s���~�T��C�S�2m
?�¾;�Kq��+��SPm8�NMGJ�v���@��zɢir�g����
{Y�Z����R��] bmU	�gd^v��ƾ�Tt��FAa��3�� ���<�D)��B����2rE��^~=w-�w�`��X��k�J�?�-88��D�/��i��*�x`]�3�����%�w�|�o@����Kv���|���=�i��3C$���噬��<��v��{�e\v���=���R��J�B8�h��TX` p�\�`�2w6�958d��CG���B��/l��5g�4�[���mP �І�E&�D��Ҫ�N����c�$$�7�T='4t��e{\9z�(��WR��&$�D��ΟW���|f�W�Mg�@�A�X���A�O�[������U��̡�F�ȧQۨzk$I��B�#�.ـ��df]«��J�B�f�*�f}i�(�s�Q5x�m^�`F�	���߶#I5�������#���.�*�_Z��?��o��#*�ʚ`p��CÂ��H��/��R���!���X��Ƃ�e	�$��1��{�GCs�6O�0
I��#�-�6H�wx ��7�����7��j:Ա��BB�Q���w�(hI�P�10щ�����E,��Nm�AW|kGWē�Q��I�
-�T�q��^}�۶6T{Z�Ro�5�O��}��<���޻�'c�X�8f��Π�f!�7D���&���\_��a'�v'�TR��=*b�Ы��5K?u͝���Ԡa�i^^���k����t�@� 2��ۖ�D{A��Y�t��?P9�=��+5���Ѐ��H>��o氌(��qG~$Wj��_Ky;����z��/h�$\���w�S����"�c�)�K�	 _��x� l�5��̚���h�.�D���3A�zn��`9���`'��X;�j+G�peW��Dw�૦�#E_`��n��:�*FiiR=M��_��ez��S"����������e���lC��n��"@������=A�y�8 �p��Y����u#?ے�J���yN����|�����޷�K�b'�� ����b�Q���BE��/���ÓU��b���&�7�L�+�V����W_Ҹ��G�tM�1s˦:�j��=�ݒ_��,�S5�dO��̃��F���ڲ��I6BDP�I���*k�#&��^���f�� V�����W��舥ݯ�S�O7g~t�6��r	1���*e�M�WDp�|�����Y'��Q¿�I2v��iR��P�O������5�g�/�Y�W�1�,�E���$}��V�s@�{�v^`����*�i$�<�@M�{%��VQO��������oYI��]�?m���f�h�� ��%%i�,A�F�xǊ�_@�+�p�j�4�]k�J��j����G�^�{�R���^:����%���zA�����>"N`&(RF��v��X�k�� �,���܋����R��A����#��*��H9kmF��O�s �%��Q}�k[�O�qć�,c�t���q��E���@#����j��0l{/cʔl��o��^�lgJZ�ޏ����3�H�'f'o���F���3Jg��W��ҹ�Ss}I��KLxXe0Zr(�C��R���Mv���LO91	6�G���n����pD �t0gi��'����I8�q������0E~9��/�+ 	�������l�����}�����d�E�N�� !/��Qe<�Y���>3��nӼ���[P�r�<�<�7�e�B�*��.o×y�G���r#�H�/ �_�l�oF�����+J�%�{V�Ѧ�W&y�hfh��EZ.XEKd���?\�P�!��A�!9��P�g͋.�ܳ��<y�4f$պ"��t ��M��-ص���T41Wr�b{v5��Wt��LE�����o�1బe\��]�C��\-�v�7�|,���]*��p������A��Q�z&p#G�d�X� �p�A�}�Ϟ�����]�RGS�iA���楸}��y,��/�l����Tn�zm� �����v�bO	�#�5�,�&w�Q�]VZ�5�{�0t#z����>�m��.,ro=ꡟP���5߁Ŗ�s��~����Rϻ�ko8$v;�]T`�Uv�W[!Jh[$t��k�3��8g�gx�'l<
W����Ĺ��N`�!�cl�P�����^�1�	K�������a�^�c���Xcj�|{0�����R���I���`�J�,��e����֢�}noA�0���Aoj��ƌ�a�n�U�c4b�.=?C�mOʙ.����֐%{=�����q�����0�ܪw�u�?�%��%_	��fq��t˷O#l%T���٤HĒv���E��^񽖚�e.S^�o/y$.���ڦ��Qͧ�iY�GI�x�j����f��5L���q��X���N^�^ta���J�d��3+^dƻŰD�K[(o��E�7E~��R����l�����v�`�ƺ�X�!(+]κ��5����d�&��KGj�~���^ھ.�(������{+�cv/-@�Q��.�ݠҵ���G��]��H1ٱ�)ș�S?�}|��Im� ��G��X�Ie0`բ?,4��A$����v�;׸�q)V�,؉`V)2����xG���V|��^f�|��|��\����1`?�BC5���s��`���87�-+�/e6�V@{�D�����N�E񃗉X�H�$�1G%�(XU���`�:�>����Q�0M �tD%l���.��r�E �X�Q�(�
͍g���|hqG�0d��u��&�N�p͇���0X�����#��sW�wU ������	O��V��6�%�!~C����;@����̷u� :�EQ�##�>��r���ҨA^����?�7��ޏ/�gS�_�9`6`�L�nþ��5Z�*�ģK @x$�����U�D�2��,W��,��n�r�H֦��fUrI�J��T*�"�yS�"�S���ԥ������0��������cg^:�����S,
���I�J���X��(O>�)���!ՁV�@Nhn���~f�ā^m�D��s�o��ܽ�T�Ly���y�~*U%�W�(��P�������);��Q�]�dY<Ef��1���@'p <_�L���z�P0k�]��f��b���EEh���n'7�	�f�n���0:�|e���*8���"�_9�ū��	6�{ 5q���r������ Ռ>��llQ��`�O�3婂��`S2��3۹�9z�������U0_��t8�-3���� ��6Y\�m�-*=|�fL@�����Sw(�O�� �����;�x_���`J�/�Kr�W�b���,J���ݦ/��2�N:�ͻ��������$V��D�U��|N�p+��_廣��bmm�j�η��Sq_�R���3Е]L}Q�����T��E��&"Џ]5�KzjI2�<D��Yt��&�2j��Wy⌫U��Aߍ,��&8ݪ�u�c�m֊�|
�\9Q������5@��5�..2C>���d�����1�m&�tU�AE�Y~��%����w�R��J�E�J}ص��Z׭��m&�X���-�����$���)�*UB��0�US[���p��
눆�z�>��xKX(��w�2��=�d
��y�����_�����Hz�J<�wc��z&v�hr����p�� %�^CL��t9x�0�L3�\[@��L(��o>�XjW[;���Z{IT �z�^����M4��H�S��|�=Y��3,
���/[��/���`�1VYE�6h��d?���T��6�x�E��5�f4q�sit��sFG@>nM������bt��:�?��@�[�qu ���P�g�YW$�`��>�2N�Q�q�F��W��A��tғ+4�V�W�h��v�2����Co,rWF��(\�H�}O	�c�h�e���+���.���ߴ��Q{!��u�/Y��eDԓ�M���d�͡�ɻ@��� ��������IT��x�=��m�3�0y�HO�>f���`��Ο�]�]�	�M���o��5%����AA�Fˁ�B��v��ÅD7�`5�{�Q��p�	!�LBp}�@�xܩ��T�rż�����(\��(��9�K˻��sY(}s;
�C��Y�옭�SX��_���ŀXWn�M����F��yf�=P���m��N�a��̖��� �B��Ƴ���Ӽ���KÖ�1�]*ey�pĻ-��)-J��h�)r�_~|��)po8K���jC�GL+�Z�<�r`a�t�8E_��Q��D-:n��A%����YK��a>H�xo���M�v'�V���:G��Q��$��|�Gaρz��;p�{���t�'�	�`�9�\��,��0�σ��݋i���.��y��ǝ:�g!j��׾Lʫ�����_�-#'ܴ�+6�%�د�:]d�ԫ�9T���.��
!��F�ntB����LS���!�'�1�_�y��ܻl�,��BZ��d|Iج:�Y�u��ǉ�T��Yf���(�����-���ѱ�׌d[���(0,؛>dr�Ym�:��NY�H8�5C%��q����[����n���Wr��of̌D���0b��N*+'���ߢ���T�5r�y$���D�~}CO=�Ĭ
�6a�JI=�-,`&��:�d�8�z��{R�:6���r�/wh�������S�J��`^,%��^.�?�NR�P���B,������V3��9�ū:���2G����U��|�g)�1\=���u�*:z߼�F�m'K-��z�����Q�1i�,Jٸ��7c^�ӳh��)Ǖ��W榫�*|��pj�Q����K6�p@frhs�}f�@Z�M��ܬ��S�)tD~Q��گ���@���H��g�Q����m������}u�,���#��ª��﯈��n�Se��j�8EN�H���5.J{��Oe��s���K�� pS����E��:;
{����L�Ku��s5!�;!@1��?��Bb�������(?���C󍢳^��)����~b2hJ&:���-V�i��R�]Y�����Je�;�H����W�B�����ꄿ��X������lr�%/[�����.��|?o�d[+�*�bӜ��=S�id���A�C�PU{�ѿ�b7�[�%j��|��J�'#+��se�ִ$GN��0��A����!�>����v���3��&��R���t*ٳx����f.JM_���8Z�@�"��f9�����C�m��?m-e�g�q>���\�8m�}]���g���������IA[��+��8�X��U�H�\bO@�(���]!i����a��"�5eXr�K�d��1�R��6~��K5��o�=�iY��$>:�:cn���3RZq��1ױb8=}v�g�/�X|7ة�i� �-�;�j}�UϤ�ZK��:��(��M�Zu��V�O�%�܄t�Ȼ�\�Q�&��׸�9�� ���:m��#�9E��*��u@�_��U	O1В7��S���lh_��%
5���x,�� �E!C��m��	<�b��<�%�vl#��d�;��Bv��n|���o�dJ�X�Ff�O$o��~����$�42���Ǟ��ީ�O�<C/�B��ƞӹ��J(٤��|)�Z�*rm\���`��q�B��ԣ! 0�'���;�9Bj,u�����8���iP���g�2��VŖ���f��9|�B���8�qiV��������vl�:^�>�=����� '�]϶�e�#~�u
Mo}-�cL���|����]��2dg%����v3�����#o�zƯ��	D�Si��a�Xj-�@�E��P����I���:eB�W��=fe^�i@�M̪��R��*1C�;��#0D�T��+��ŦT\����b��ʍ:&O�3}Ӌ�H{lʛj���_�	�WW0�%���.-WVUt�>#fp|c��URy7H^�hA|
�!��"���g<��YY ��i{[���;�����.$�#�H�u��k����ǘa�.���ŌY��yb�<�"�<`R�cɇ'˙�Z�zGwO{���wCođ�
�k��Ѳچ�L`�G���x�.�$������Hm��7�㼮P~��1+�	��v|c/�>Om]t���7��pۗD�͢�������٪{RnD_�rȰ0JG^�;��_j�����o��הn��51�荍��7^"(�56!UF��u��?ݗ��V;�@��_��1ƭ-x�]3e��hʵ�����O�@i�DmQ&�?����u�gyta��3�Ӟ��o��km����jE7�鿋\���+�&�1���Y��U��}����k�����k�vN(y��\[�3��pz,����)�O*wx��}qE<���H�r�n��ј�^7�~&XL�~�\��[�����l�X�?2�ؚ��W�)̓���6�V�p�S�vl��=���f�d���sb�Oo��mEl����h�$�u�� ����N����W��τ��G�ͥ�)�ٽ�d�_�����5��2����۬��v��O�0��l�k��'�Z��l6��`��7�s�:�F,z�z�oZ�[�ѵ��X��[���������i�3�w��N:�H���è��4RΘ����e�Ԝ���f�~�kjz`W�/R�S>�S������
�#�1q�8�g��,j��'�PI�_ �]!�S�6A��>w`1�C��� �\��{��%B%�@����J ���Q^�9�I��QN�%l�9�Y�<IeM��f&���C׮�Ý���7HO3O�!lN�|�4�0y7j�j!Cl���c�aJ�����%��: 6 �1M�@(�賁\X�vu�2G��0�F�������ys��Q��MXX�m0��i���b�z>�>$��z��ӯkj�j�̓o�!��0���x\��E;SZz�)ϙ�t�~.㱌�4���*F�L��h��蛩n�u�KH��[?0��� �ȅ�����seŜ����g�ז�B�OZ�8�_����1���xp�?��j!(8?�%9��B���/2^�rE�Y��)�������	���r.�]cf\aG���\=ر[�:�}�H�Liţ������\z�fmZ%�� ZӃ5�5��!�N�N��M��O��W
F�6�G7I�7MHJ����;^�5Rߕ���s��Q�6{ho�]��2��BE<Ɉi��wRV��t���	1��fU�L�I�1����/����#E6���s߉�Ѡi���@\+�ڒ�4�H��x��L֌I�� /g��@PP���O�Mv�H:�K����)/fZ2��@��3-$!Jr��xh��:�?��#�����|z��P�7:���GD)�(�V�B$��#��Q��B!@~Ԅ��7��[�M>�kw���I�)ɭ&���l�:d��.�Ϊ�eѺ�ien�3�&�\�X�*��q��K�\Bc�y��� �of�Cl$�"2��s�8�|�Ps��ƥ��X>x��C79��j���萦s�8j�m���pDp�F?��<�B@�\�Fov���,�?����FVjɴ3ת��[��c������������,+�*S�Mj��K|���~�2j�a����k���Pϩ�F4vN|�
w�����N7��w%�K�ut�-P�t�W�������yA͢�f������jT��g2����l$�X�V@/˔�:�X~L׋�j��`������@æ=�l�>�Է�޼���Ak����L���3����V j� d����=�i`�
D��%r%C��;=vw�uڧ�Ū�1�nPIe�,�s���r����p���IQ��橁 ��$�7���7f �Y֪��b�<�(���oM}�*o�o�m�L��0R����I*��XdqBr�A�X~VJ��Y�C);ة�n�v�eʤ#�k!Iv&X%��d�pj
���UT:���]��N$�D�=v�'�BѶ�3��(��܏S�n�P�:e�@��~c<��\|��i�o�f�)wV��XX���X���\��m��m.7��]����E(�(C�ܝ]�&RB�=Z_e`��H��	/?�������)(��nU#!����V� a��tyZH��x�M����>���>�=&H5zA�0��e�T� �`�|�-��d�� g���΂z͞��WO�����:7,�!���ʸad�̉s6Z�}[�źv�Yf(6����A�/����������Kip��ԑ�w�C�ЃCC瑡��I��*3�誳
W�d��4^�x6�;��	Є�p��'|:�cF��G����LD����x��Wgw_�O�`(�f�X��?R�*��� �L���y��9�V�����a ��`5)-��-�՛BL���Jrʏ�x���8n�p).�B���'&\�O6LDj+����:M��8@{�>/��NO�V.�jrZaQ֥%�4�4 q��	)-��H�W@wb-ךYِY����g-�|�l�G1��zE��ǰA�YE��-a���X��+��A8w$��C������Y��|V)2�cO��>|/;��\?��?{�:#��+�՟os Ӈ[D$����M�1��(�C�����	z7�x�Wa�3�C�/%d��h�``j'��KG��~���[;��̤�_��u���Z?[���q����a׉U���,�W�\�}9�b��>ц�a4�o�(\dh\����9��|�55�s�Q=@?��)Z��_
,9��9�����B�}�D=m]�,�'���O��v���A���]�
} ���9�us�73�V�t��4��%��B��Dd�}�����֒�%wxP\�wb!����/�u�	 ��H�����tA��������N�����7��N�H�#�lmC:�|���7E�����QD�ߘ)����S�V[ɂ�U��-�c��
2�X_�\��A��_�[��<��I^D�CXp��CR��.�5Z��5�����J���x��#�`v����^�WY�4
`����+˞��$4o66�Z>x1iVMɣ��I����X�@)��Bk�+���LTxj�uW|�C�:�5Tք>Tu��C�թ��V�&[lҭ9�����U�t��X� ����g�9�I2�;�0ɨD�͊���N���E�V Cvp�����̧M���<�u$�[�1n�N�g�ĉ	X��l��d�uP���w}�K��M�o����:��
����d�H��?V%�����gP���T��A��2�}�-�hvW�Xa{��k�Ұԥ��?xraX�Ā�>c��K�-�(؋*Kˍ��p�C=k*7�}㝈��Ζ���lH�dbV�_ۄy�V,�0�$�-�S�4ޅ�j�Ț~�� �	T֜[-JoF���n����X��R�粋[�p�m�~��A�
!Q�����n�B\vT�ӗhI�4��5�&��wp~SXe�׾�5X���9�����M�>i�r��_�Ec(�urr�V��H�s@��?��a��1�AZ��q�x$�d��˧�#�>"��AXE��RS��+�D�gIV}wOx�/_����/�{Z3���{�铢��~�2kua`��jd���!������`����}��p+��0,O��H�W6�k�������1E��k�(�+K�?2�g�V��a�[��~ZR���b"��L�'Q�9<�L���Wv�%z.��݌U�	=	�����ϡ�l���[8HU;�)S�������g�O���
��E��D����m�.���4e+0i���H�ۨ1N��_��{�D>^�W0mm~�B�]�m�m�]�)~ƪBq]=�k�k�G��9_g{���q�tc�e�f��[1�����h/�i��o^�! ���T���u8 �n�?^�uy��ǲ?��2nҨ�E�Z��d����9K�\����c���� ��$��_c|#iI9�5M\aD�?]	�N�-������(�^l����5���H��/�se2�n%�h&����b��!c����n��
������_�^�o���������S�鹀���
�buk��&Џ9U#q%���,6�n�E�Í��%�M���'J���^X�LC����jP�	�R:�P4M�$��͘���.{Aֹ����>��b�h�_X<�@�6� 77��մ��ZL�z�j�v,����-�ۖ�ccM�ӏ��T�	�� /�ȳ ̔��d�
��W����J|m�Η�ַ��M	����,i�un1T�#I�Neojx:=`�_��Jۑ$�y(�"s�$���C����[������\b��A��:��V�H,�M����V��cw y���w���)����EK��5��"�Ց�Ӷ��NN��e�N��Pq�%��9�\m��R���&��^3�_ٮ��P֕o:��*�����|��<[�gt,`��{n�Q6��[y�6|<�	�<��(��<���/���E��%_���ٝ��˝�#Z��g��:��q���(|��-���o��u[v��4V�Vh��X�cj��y }i%��%l韽�*��c���2��t�����̨��qW�e�b�D�m����*p��P�D^m]U;"������d��7[lMl���>��þ]mZN|k�,՛�*}��4U��'$/��X]<�븪{��*�?�P!�;���7~I�^|�.@�� &�Tq�\��8�k%ɂj�>�C�vS�jF�Ngӓ���7rQ_�nmQ�mA����8��g�ې�ͯ_j|������#�^�&|$�To1��Mg��X6�ɾ��0�N-����|�b@XoM�'i1^���+�!~"��~b%��VLi�o��-rK|
�d&�S�j��������sv��\�����cM�G4��OGX���G�B��W��p��XD4�L�	�~��hC�Z�&��]'�5���)���w�?��Νy2�މ���z��x��a�W�Ý�
�����d�##��������Cs���K�o�~��[���osL! ԏX��+C�tB�.X辇��oͳ �Q�'6�}h�o����e7�"G�W�Ӫ���j�L.o`*���/\>п��6|e�M�aȎa%�>r�=̍n]�W�'w{�?�x�\���3[=(�_�4�Z���q�#�� ������}H��3&/.Z|�^3n���aM*G	~�-'z�3J�dؔ�����a���I��g�;&m)"徻��6e�+?FZ>�j�fW9Cݧ,F�����"���X$��i���[�ĪZ�iʥ��c��G��_��T_^P�h���)յ��O{E��ؔ�(�*"x�0���.��QqE��p�k�l��ѱm�����+Z�������K��땒v�V�������.ƚ��_�ˤ�I
H�c�[KϬL�w���
_�&�+INC�< �Q�ȥ�R~���#�H?����M�GQ!���*3:5=2i���0�I2�
����6���mc��tKf�RiJa�Ut�G^�][����/���rs��}�RA����[i2�2&Oz% ��Zjŋ��O���2�x@Xr��+����#wHv�B��8�NE9gye	|�	 B��ٱW������st!�� �$�'�뜒w����qsy��	\����!����?Hlbn,�qу"��&.����S/�r���s据�e�.GqVj�t�p�Lb��t���Md�H�?��i�;��6s�P"�<l�I��6|-���[���� j^���e�n��NH���P���YYGﺰa?�g�많�FI6�)ҖT���[�ߪ��S�U�'ض����m��U�Er��v#�O1��'\�|魇�u\�̂L����u�`�)��X��A��L�#\��Q�n"��DZ������ sm���);�.���9ݿG~N�k���c~���P�Y~�)���?\�oU��˄�x��l����n��㻝It.~=�4wm�Zz�R�?����.?��%~a���/�t��⮔*���Z 1�|z>D�5�[�?b7�e��{�W����#��K��r�2��*w1�8(v����v@���&j��a� ����)�o����X���?ݪ�v�;��+��R]��'Q�/�N��[sC�~�ӄ�E9y@H$�}U�XFg$:
�cO�%ڈ��w��b��DP\���R�ݡ��(��mm���I|�.;�!��aB��	�{�F��<��ο�<g��{���GU�H(�7���:d�B�0�:kA�]*�ڦ��r� j2�G�v�D��C�dPiu�y�H��(Z)ɮC7���RW�u�k�m��-��Sh��#�P��(G݊�X���hz[0��{����
��!�}E��_��4Fg�9��_�@SC6���
6��D��Atͺ��0ח!>t�b��O'�`e�<[%Um��m�;:�l�Ά'���m���g�3����r����|����G�����P9xQ�b����R���o�i 鈴�d���SލEI���ֺq��y�2x�*weo2�p�I�aG�Pk�p�;ܹ	������.�j��ޢ��n��)���]ͦf�_�@�2'Tag�l@����zwJ�cX�a����ԑ�ߌӢ� �|�����G*�d֠��ˑ���8=e>���M�S�!h�����8�����ʀ&@z���*Mu�i�V8`�Yѕ�[Y�7:�.�ٟꌘ�x�p@8g��>n�/5ie��NF�Eޔ��o�8����n)��h�	�8a�l(�|m��$��	����h�� ���78���\h�),_H��l������j�6"�k����2�$�^E?UO,c\��d��QW	�x�-�0��ЅG���u�a�2��;�*g��hE��*[�.⺪ǣ �@P�k��2����S�?��ΰRp}�[�Q�����t�f���#n�����M���͵��������G�/���Z�C�`=�=��y��¡�R�t<�I;�r�jXa��2���lK�^�X�,
��!�)�.!��yT$�/���)��s��|���)�\�u��M��:!�������	�u-����@�� bH���X��rQ��N��:Ae~_V"?���S	�:��r�lϓ0C䄭�a�ؘP���V�n�0�]����%������2W"�2l�NAD�C�F,��*_D�_@�Y Fi� ���6hF/�&%��&}��Q�y:�-��I)���E�p��͸�D���[v��ٔ����4X���}�HcC{�������"�6�	ڒV��7��^��*Oo�B��k֛/�f��e.��z��h���������P<�b5��`(���z�c��ZZ� �H��է6-)n��]޶��/���ûO6�y��z8n#�ڇ���2�u^��h�O`�b�lJXΔwXQ�Ut�b'��RZ����d���1Fߛ��S�d,+����6@*1Eʸsb�#=�U���z���ѓ��� ��BN�2�z7�6D����e�
�k�뛤Q���E�wΔ{�Vq�a�|2��6�5ڌ�W8fޝ>I��]��bC�{ ��M���*�(����'�iG׌٪	ցK��{{���c�n�t�+k(��ϸ%��`
�$�K��T&iB)%NM,(*���U��
��#]%9E�Q�Cv��l5c���˙��r�v�����
��wF�~%��W*(կ�}��_:#F��x�xk{�J�~�·z}�U��П����d=�17�H��2��It`ۭ����W�> �8�á�����-f��Z�׊�/�v{� Æΰs�}P;EG�s���VU���+d��tŊA�fXV���<�0E�B9{:6ͻ8�x�������`�W����ul��e�kǖ�AoIDJQkP�cRդ+*�%�ݗPL� Ι[=����O�0OII�x��y����E������r��=����N|�#��?A�y��1�Y���L��}
̛B��|l�|{�������zg��@	����v��3~�B�L�h��CMlM�yS�H'͡�%�k�qx�1�l^��0ݶ6á�X��tw����%j"�8�X�ԟ�����;��B���~S���X4�%hX �Zo��@J�u$)�֓4��ם�x�b``4tÐ��ԧ�>�7��ú�dǪ�	2�se��k��)���������/�fl�}PYx&����œ!�?%�9{d�&��w3J�C��J`�j��u������x�: �	�洊�W����@������/R����Cȶt��
�೽���V�$�*��Pk�}�&Oc����y����e�3CC����
S��X�/���N��/��ef�)o%c��I���,A�F�sц%)�I���lR� FY;n���ޏ^V��;�d=��r��E�Y� ���Pe�5\�Cq(H��J����$s:�J �7q��]�˚�2l�o��=�� �pC�H��{��[�h�`<� �&��Li �뚔��P���]�.O-W`.AN�ouW�O�;��)��tDǩR��M*CQ#��@�����!�!M�1(��	m�~�L���f�a��x��r �Y��Aݧi�G�$����ɿ���Z-(��O$y_t����Z4�26���ǥ��<7;�^�n����.�!��V\P���'�b�r�[�N�|���Y��X��C&�F��{6P����J��ĩ��fB"�~�I�~�l��N�B,��yI����%�w_��?��r�Kᯀ������J1ˋz���6#T��"��n1�pi�"k\�.&\-`��&���~^M��Ff��܂��_���O�W�2�_�	�sM���b�9�_��uM�{��5��C!�wcHA,���i�nC��4�䫧0��}6�ǐ����*O��, �n_��m
����W���$iB�,�$�:���3_�$���^]]���T7C�m.�g�e^�e���L��<_���E����YIa���Fs�3��&����j3�qxS#_�&s�R��b��%�x�Xؒ��4�d��>[O(�dŁ�ѿ8]�������pT��Mp�J�򮰨"��\Z�s`�߫+��Mn���T�aU��t�d��k
��:$٥ٺ�4���'��rTN����$le���ms������5�pw�]X�X���^et:3�`|���Ō�2���5�MtN���7������X@�7�7[[��j[�5F�H�~C���D;'RF�S��p+�X>�<Q�83n�ߊ ĩ����Z�Z��|��q�j3����2�+��������h�Q��c� �� �����O*y���r3)1W]b�{��z=�}J +Ʃ�PG�i`;\�h}Am7,����� �Z�G��]�vXG�R��������v0=#�@��.c��Pk3�9l��;�
�4���hR�*Z<^c��D�~�m�AE�T����ʯ?�F��D�zG��$��r��+{���EOn�>��z���S�~*���w3�aR���������/jns�~x���haՒR��?��*�]N�͘n�$+�� Cу��s��K�.±O���r��S�gg@���w0���]�LN�,~�H�1���8�G0�R�!H���a�k�������q+��$u.'��U�XR�����-�*����~��'h����w(�������n@n�ݪ;��/�& �ތ<����z�쾱x���"�B������f��R�������21�PN���h=b|Pekph���;3��+��cb�!�B�1	�mr���ض���l����k�/��BY/E��5�1<�3��]vD�{�LR}��VqI�1�
���,����M�B�?�ޚ�:҉|p���X��`Em�CXa[���z��w���6�%Sp]I�*\�~�E�����i(Q�J�;���/+HX�k�6�:�X�*4���?��I5h;B�۷r���2w��J��#M�>�grt�¿�P ���2��=�0�b��"��(�&����t?���`���+>�$�y�ٮpk��Kk�L�o���ЯD"s��	��=����0�35f3/�Q֕��	0���ӯU���dS���	5.9�����LrFk}%�A��=uJ�'�pvu�?�2.�&��(��3�L����y@����r&�ƼQ��rZV���+ؖt��n�����T<Z>�S  `2��޿���ZQ�\�N������MF-�	�%G@���ư_���Ӗ��o���z�<E^�+���!��E��C� �q�.�HnRH��O~G�S�`����
��E�W���Σ�����W���^����Cc�13�'�YU��Т�#Cȴ;SE�F�x�W��&3�:��ԇe��pj:���1�����ȯY�%jZ��ꈴ���m�rG+�~��)`2K���u%,b~sCi�~_���!)��m�ة�|�1����qfe�{����H}�A��۔�o��9�ai�f�ѱ�sD�#.�ނQ�&}�*������r���tbx�3i��^�a�;��4Qls����+�-�`��[�98��Clb��B_��$(F��T���oŇڂ�YDݱ"]u%(Iu��,f� ��w�H9��~���)]���[�;������-�Q��֦��,xnE�0M�	�蜙����0��َ�)���o�]iA�i5W�V�%�Y��x�D@ķ��0�B�vY�9l$vm �&��Q�Ƨ�$/�WT��e%D�_� ׶���E�k ��|P[J�b\��Ę�}�ui)>�*k�#T"\:%�`(>���s�Od��cM�1�>L��	�ĒJI�PUd$Q,}�)�G��]äV��\sBPB��~t[˺ ۧ�(�|޽��԰�0e���"5�a��䋁n���	0�SԉC�L��Ѿ�[��7��Č�'3�&Ô[�M�>tu	��t�Y�6wz�b�Ç;�g�v3��x1uW#�9w�. �2uz9�MH�yz�ϐ	�{q/�P�_��2]��}�꿍# �{_ɰ��l�C�hy5�y�-�1[�I��dM]<�8��a}���;��Q�:
��`���9�)CmZ����ڦ}:�����mQ�jn_;lԵ��o3�YY)p.<1�xW獭���k���~�S��>� �8����������xo�ʉC�c����K@�O �j]__NL ��t���E=���̱C�pW����6;�yw h������M�I���^W����(��ƊӃ2�7hԚ;P�C��EY7����+L-V���^�~�J�}7,���W�G��o���B��hQ�rs/+`k�1����m��Ը|�Q�ؐ�-������nv �"�d��gX�gk'��0�t�ňh�[זD�[���ld!���\l�k�o�ۛ��^���g�ͧ#�q<�oI3��l�U_ߑ����N���3G�d�I���C����@��vZ��I/���؞�������$�J�\ٞ�	�"��-h���_��$�X���2���k�T�H�]$�Pֺ����Uf���w��o���@c3Ku%p�FݛA�h?@��z;�ϳ���}�̜�����w��*�h�Bi`q���ʢJ���y&~ڟ�t;��_��d����})��#@���%��������,7����z������,	�<��|�G�T�6t�^Z����\�cWW8�p~�C��Wo��{<���{�����A�[W}y�su���Gԙ�h�'�O�r�$���ຨ���ϱF@(���ۘ�	ڸ�f�scxQ9O��%�36�lxB�/���[M���ds2r9�0�ҧ�f���7��CZ-'أr2>Cud�R&���я�
��V9��V���t>bV�.��yTڎf��b3�׵�m����R��g�=�P{�x��Y�Ж�H�.�~����%O����mO�&�T��z��3a�%�BT��+F[{�!�ۜ��.��n"�w�o�깝�Z�z�cY�<��f�+���tڙG^3��+A���z�]a�m4WD&�S�D��R=���׾���PSl�U�����,kH�$�	\��X?����T˂��=�����7�3�Ad��ǒ���d� v�*8=��[�8F���5m�s��;�۞8��O�K��<�x���Ɂj�;i9�c{Ha�@���3�='\e���\����/"[p��-�2^��0<@s�XߕOv�Fp�Q�]V?t�s�Cl�M��4�b}���(֟�l��!�>��9Ё��;b����C@�tW�[c�]<]䫊�wN�%$ɯF���u��6-����o��@v������ڀ�/fF������UV�������	a�el�̟��� �g�{��p�2�}rI�F�z��;D~�^��`v��5ޓ��=U�(b�w�r���8l$3?3��~�0�J�%�yg�N�=�Uկ���^2�PԆ�!�v �)k��u$Q�=C����i�4�`�)iT+��L�����ֿ��s,����l�b��r�nft��u'h����x-�[-"|Q	i�~)�8�խ��𴂸�t��bjA��YG��3Q�n�L�8���N�Q�����H���Es��P��]������8�v(��q<h3S�0h��O�X�O�v-tf��[���kӅ�%��7�í���wN���e��]��1�
�XȨ)�w�3H2J��&�(v��Dwt�ͭ˥÷0��ޘp��ӵx�0�%qj؛��^R��Hf����*#ͳ��8a ��h��"kWȥ��ч嵫<}�H�9����ɭE�.�t}�&NC�
�n�l��������70ǔ���,}����Tg%�6=���<�E��w0�Z[8T��b&
U�a�M��jw߅���W��B�+&��l[�LWP{���Ĝ3�
�3��P'w+1�7c!�	��Sok��B{`�7���ѵ2{�g���!̀��a�7\!~��Ύ����T��-���N�gv3�_��#����������7���?��k�}{�8�d����I�Km���$ ����'[�
��P���L��K�^A�p��-��b��>ӊ�-K}�#K`?��zF�f���51��h�Kv
=K����L���ǹ��x��V]EA^X��{T��Y�E2�
���¤O�!$�L��p�p��ܓ��,�]�Dp��d?�����h]ۦ;�[��Z�`9Vȕ֢��j�c
�a��^,��+�5T��s�N��AK�� �GG �iC��S�h����&a,�����m�����t���%E���Bk��N��Զ�ؤ���3>F�F����`�3L��̤~VnL��`��C�j� �x����V���&�� ��e���ƕ�p\kN�AwVdDK�6��6�[�h���ܠ��x�#oS �F;>^eț�a�,dlƳ�xL�9h���l�Q��
���s 􄹛���Yg�������ÏÀ#:��,��k/>��К>yB���l���oj -"vz$He��䆱آ�=�Uw��M��h���Z�����A-�@8�s#�_b��������N�I^�Vg��A�/�]Τ�v�.�QڌtN��5�����G�$p��m�I��~��~����1��h���[�k�7ո7J�q�%_$X-Yj2?c�R���	F��m4Mտs����^���5-4ipu2�јY6S}k]n7D:�!���;u��\̛���G����<u0���J�$W*EtiJC���,��^I<l5�5b����Zk�C�"?��ip��/�)o}J�cxV/���ċ������T�*t+�[����3t���H���f�	�漬�*�Z�	���0&Y{"u{��1KN1ۼ7����"����U%@um���+��3�S��6��L�CɏµR���^{�e86�����a��ɰj'@r�� �����ρwUͭY�&�,v��-g;��}��0؉|��݈�!p�t�2O���o�b�9L.Ӈa)����u�x|�#\�����r7�4]�l��ү4�,�l��V{"V{�Y`��U�ɿ�\��e��"�f������5n�9��f}�w{w�=�8vVֿ��h�Il���L�Oеe>G��>�;u�p�|�^���G�>�}�P�2}x����o��w�q��J@:]�w����	�=���{t/��	bm���.�j#�6-�
�Ȅ��卍\>(�hi �D��Fh4�-U������mg��ٱ�^J	V��@d��l,2S���ۡFa��r�����7����1��d�hmCH���{��a�aJ���G����m$&��0�y/�_�g�q��J�2���Q���M׌�}u���dY%!���%��V}c����ϧ^���\jg�t|~��!�[F��4���^Wb�vc������z���ۿ�����K�00/%����E�j�h�����ee�*U���ɓ㳳<�I$�I��k"[��}�a�5��d5��ԫ|�o?,?�2�����y �TP�rv�;�Y�#W>�KDZs6��]Oʄ�����5�ҵ�X8�>8���)W�m����c����|%L�X��O��^]&�,�׊��0ZD3.�
���B�*Q<ר�.T�nq�c���9��Cp1��S�(�L΢]���]AT�B;�Ώ��6e��]�J��܁B����d�� ��� K�AؘE�
W�qb{�Q1gS�9��
+��ph�<.�t�r�f��O6�.8�	���|��E@�_�5g�輗ע��MPlF���lF#�l��g����څ%���/>��,��{�SN�`�*�VX�2b��X�(bc>̒��S@J���P��w�ι]Q�3(g#��oyǣo�E�k��]�#�9ו�7���G�w�wx�����>��c&A�ޢ^ƭ��J,NZ;��0�%��҉�qa4_�ŬR��Յ��̃�#�ID���(�rëM"��ϊ!�0��`-��Lѝ�S���3`����]x�~���9=Uqn��ڲ�@pC�+�`�7镍z��mqt����Mt�`d�H����z�V�	�T?ri��e�|i�5�1��-2�D�K��t� ��O�����|�-��#�Uա>S��$8[M<�l���KH �ԛ\��'��AӿyF/  ��3,3�L����wf�و�7a'n0�vj�6���s8WL��R{Yc��a[=���pnsQ���p�?�"�K8����gV6��sӛ=��rE���j�I��9"��!տ$�u�҆�Mi�d��#K���"<��{1������V�T9����d�ix>5^?Έеt��E���;�ϕ���1���; �{������i��s������M\/�&� �D���q�>��%q�^�vZq��I��|��#O�;��f��D6�xT/z�G��c/;�H���48�f#(��� �(���G\%1�p4l8^���k:��ќy�T�	�LQ�WH�c^� ��wM\+�d1)�Idl��8�"�3��<�9��^�sxI����jbd�O���Lx
)��w�$aA`_���!k����=��V��<�o�	B2�'��@��˿������8��ݴwr;�)=�Y�T�$�hE��:۰e*n3_X�w�@�W�dv�v%�,pX�o�Ѽӣ�c��qAD�)�	��7W丣��4IX���lP<�������X{|ߓ�1� � _Ԏ1�~�A���L�Ye(Wc[8�!;���^�OlA�rU)�3W11U���}�f������5��i�����MM�W3��ww�J,� ��-��s�5u�%�3�?�>)HG3�)� �x@��9�������o�~��η��y W��A�*'n,��F�L�aR�J�{�7�(��+��z�~��*�ͩ�F��B�(0�"��/�M�b��Ǻ� ��&�(���x̓|Yu��B&W���ئ�1HmO4�����;P���鎝�}���ȿ@�|~z�%��G);��f����� �tg���H�?Z��^�z��q�=��5���[�(<B�ccH*���Bv�nb	������������N�J��~��P8��⣛�;���S�u={�NS���:����|	�'�7��fy:r8�����K�g��Bj���y�й.������%:�z��Z��KG�i��q;ww;wQ'�a �#B���В��V��o�l����	2���@��nq<�kP��&e=�H'eJAWΜx�	��d%�����[Mi�^W~����%�'�%V�t���]�"KJ��|55h�qGжS�(�g' ��r�. �?��f�������iƪd9�B�:)�-�����jJ1�H�o-R��p!��:�8�,�G@q��ٴ�^4���T���`��q</��%Nǽ�m �Ͱm�A/8̕+�� �UuA0QΓ�hVk����.��&��{�pVw0�W�6�B>U_ܰ�ֿ7�w�E�>�"kųc�>��ש��Ŕ�)S�"�!.�GZB[�=�\���s]�B31R(^�Ş��V��x}�z:qXB ��'$HGA��5��<���ea<0���zA�D~!n7	�-Pu�� 6� u�9�n��^�M��P���������5�n���6��I1��5��g{�6�V��u��"x��W٫0���h�s"賮�E"J��CM.�Θ��6;̶g��B'@<{&���g�&��I �*�} ��6������ӡ��E�����u�q��M��$�����-:(D���M�[C8�#�*�CFc���"�+��1	�x]Or� o
���Y��"ǇA�F�?7S�s������O����L�-�:H�Z�ӂ�G0� Y���X �0" E�>#��kG�ȇ���F�|��_P!��+�ӛ+���Yk�z����w�F�$3qc������Yǹ�2w�GQ�\Nq�`�,!Y�������ƕGO���^��CZ�8FVA�5����L���5=�@~�>���&�S5|��o��9Q�â��#'^淇6:�0OR�t@+v���q�k�N|Q ���1��h�/}t��$��D�3D����S�=sz���	��b�uh�����E0�7�ߎZz���T �>���1��C�z5c��&�����)��%��A>B�ˣ�,l��
ڸ�{�IՊ<�����e��{����u*�,b0>�P�ɥ�����&�iRĠ�e��Cڕ�3Klr�����얛M����mC���<c��4�sTpBG�y����?	Q�ٱ�l �����I�w�����U�~��;Ѩu@���i�y�4s_�CDE�VeeLϝ.������nd��/|yǬ�8U{;n"R^�����B���K*��y�$W9vT�n_�?D�X�	���kd�	7c2w�ǉ�:�y��u�f���OQ��#���`!z��%��C����:�����!���Z(��@���*��%�7~��M`s��j#��oXTY0^/��b��eK�^�۷��#�q
Z*�Ћ�zؿ:Ǖ�;k ��~��k�c
WE�����5\c��t�����Kv����jUʮÀX
<[�����ج��YAw6dK�@5��J19��8e�
����BV�{�)IJ���gy55�C[�.��p���!xYt�ȵz�.����_i�&h���oN�F&[ٯ����Z��C[b�`""��,2�x(X^��8��}��Q�@���'j�C�PI*+��vo���d9SE�'T���:$�8��{�O�(��"7S|�ʎ�����ǂmNC�w�`@;T�eֹx���q�'�5�+�8�Rv��<�8&��^�i�B�*R4�q��2Th����hĽ������<�g�&W�"H���x�#Ů���w�8��!y*M�2o/����i1:j�{c"�CV���@�λN���*��FU��lNM`�$�O����ѱ�]��q�E:�9�n�]����Cg�YW\��oi��U~����ߺ�����������o��%) �P#O�{��,�����|���"q2��h��� |����1�?�sR0�!�
ک(�v.�m�n�RI�v�,��(��2�$	�A��h+>da�Vļ�a��8#�kSq��)8"|:���b���r��� �t{�YV����w?�m���I�߶�y��mo��?�.!z.�{v�ɹNIV�X���&٥� �~�Je=[*w�ڇ}� }��^D_�M�R�ɞ5.	Hon��3<�F|���N��x��la�[e��Bl�B�\���BB%�u�]��/5�GkR8nn1aA�{O,�g���{ݜ*��b��?e��"�o�7�
(c!qX�c� Q<Ţgy�� ��64sn��ʈ��\0�t�a2Wϱ7�Ϯ��*�Im.�^ʳu�4��j��� ʼR ��)��atJ��ʳC^�X?������3�B����~_�h^JzT6��������5_��vc_�]�Ɲ�r�r�w�_�$@�����G*��_R����%�f�qܥp#YXR�n�>	��
�IA�g��� JB�������w5�7��,7q���j/���C]�u=Ύ�c��5t6ߜ)�@7T�qX-�`���g �y �c��L��OcZM��z ���P�Y_���Rʖ��]��6�4�kwW�<o������Q��{��B��q8U�5�j����8�5�<���ٜ��.Q0��c�
=�d�1鎶دr�tp�ܻ0�<�i��Hl�]�uM˩�P%S��뢍<$c�:ɖ�݋�2��A,vA柍5�<���B��`Y�^#�vX�~1hGN�S���#��X�"	����~��	TI�%���`ڜ��C���Y-��� MB�5*K�\�Xv~P�T:�����x�D�n�aR=��*x*&7��r:J���|UQ2�a.(���F��-�+y���7IIT���AbO�V��$�Ŧ�A�p�o�[���!�E�� �x'fh�^�����:�F?U_���Th?p]�X�;����G���S�w��z�j�͢�0�-��I_����Vfa�ٓ�����Z!Sg� e�o$�۹���g�o!��gp�	�e�A����$�
c���]s�����K{���SH`��������!�䥉���y�H�?A�`��}�������������j�i���=Ƅ2C	t*�?���Ԇ%��SWdzR��%�[���I���X~���s��ҍ�l�o�j��5ҞmS�@��k�'ք8����6�9iuRV��1)R_����Rf�{�e�?�y���\#�[W��F+@WΠH��iWg�ʠ�JKx~��i�\��p�k<������[C�O��,�^6��!#� !���J�f��[��V[��PVͧ�	}�-��O����T��0��9?|��l��e�n���`���S����(���6I���.W�]�΂}��^S�=x�E�n9��`�h5�s���B�{�����宆c#[�D	��'֐�I�)@s_��HQl��Z��9�ϬuW-��|X"f�jI�>3ǞXH]�����)�[|Hs�1`q������TD�;��D�~/��.�]��=F,�{w�kj�0{�����S��<���S^M�a0����/�)�Z�f�7�7�L��CE"=�:���H��� �M��"QxM�>�,�]G��gB�<��G%P��F,[4���C-�3H`���b�+N �t���beu-|�+J��;+4��=m'?��,D��[8A�V�z�� "A���Ži,cۿ�K���9IWĭF��Sг��F�<{`�N;*R��1!�=��z��7���b�z_�| ��O
��> �AR��-S�#f*-|�ߘǚ;�#�As�Cy�ɴ����N�?Pe],@��5���%X��`��8�z�t��ieb�H[��w�Dh\Z�853۰�Ys�p�zv�B#@��ͦ)�EH�E*@����a��P���=b�+e�H���YlxP8�O��I(�ڛ��"�r����mY	�3Z��:�����ɕצ��Nm���"�W���ԟM�u/Z��/i�ݠ�D�ñ��G@�b����c��B@���a�w�E[�g5kJfU���,|*��w!tg�y�u9��j.nH3/�/�����#�ҽ �����1J��0�k�_�E��?/������4nk������M;{��1��媖��s����������P�ق��[���[�EG�g.0�,D�D�gJ�pNKo�dBr`\4�����ԗ�G۔�޽,���?��~�%o��Id�4��yb^�ǋ%�N�7�� hix40�N�Zʶ/`5�̶�����H�v�w��1y���F�"~^`��B0�, إq��MpP)���������I���T��La�<�N�~ě�)�o9�����F�2���}÷@u`�n%�J}jX��	e�j�A����s�کa��'l���o�;�ql�`�|X��Ko�Mu���H�S�z??U{)��i��rD6.���"�[YMvn�VGL�`H=�����E^@�m�~��T4v0��g��%]k��=�d@�b(�@��	{��?��pT�(�H�42�޸��p^��^;!�q�¶f���:���������l�l*a�(�a�r	���j��y��]����h�L��A�U�(��*�sh.�/��cq����8�d��������1-�J��[��{G�r��_�{!��`Н��@�h��:-6i(���ڮ����:��X"|��rf1w���ڙ-��@8Ƌad�J\z�������dUr�'�ם��M�Ao#��+��P'���Jz΃�#kn%��T�C��&�yY���&c��4ra. 16OW�h@�~qN�M척	���d����;>9(*��}(M�2\���A71��X����c�-��y0�%`R��ص.�|&b�Su*
�sϣ� V!n��P�-j8���n�:�R�.����}]�����̧m�d��׹��80Hq�P4��z���o�mˎ++N*����@�W*�ñ��El&�B�+��:��W̝� �2v�e��8�vB�y�8��ؿ7���G�����eIrF����U���� }<�b�bb������֫�d|S���.N��~�V�c��s�y6�p��b�q��r�Fa�h��+M�q73*�ǣ.Ue����f��"���ʰ޶7�E�1
��$\Q��zWC��r:�Y�I��K��^���GG�Y��Փ�/%6� �q|/NBm��d�K���8Zl�`!ӓ���*���C�O�|xQ� Y����!d�h.6`
��B
���ӏl>!܆w`§�V�.{x�	E�Y�E'�'�D�p�)
c�!BRP�")GY��OT=~�����%xb�%>��>�d���}��n���E�/��e���z^:�;vZ�[]�e�F(B9uY8�Bn
r�j2���R���nhb����'�a�;���q�Ap&�pH���/��Ͱ
Y����i�����S���Y>fuK� ������R�|67�E���Yy
:�.0T���t���|�����s崎P)��/�J�9�29��B��.�T�����_�N�xc¹�b�|���/�o����lƥ]�K�n�d�^EI i��=V��? ��[���w���t�F+�(C��Gm�a�l��@�e������Vhrr��i��C�l��� 9M�>�Oi3�;��픫J�k��Mf,!*�օ1����T��Y �	#0���~��(�aqs\�ޟr*����u���nu���f�6J
%�?5c��S1Xv�v����Ry�'%!.>�U��!��h��B���.�nQ�mǗ�w4z@N��3��mQF�ꄳQ�Kg��h�&/S���㜚C��R����-�v�d�C15�7�L���Yr����n�,B���o[�.��)Y@�� 'SρT3o�i�a%�Q.�Bg��t/�%�H�h� |\�j����_-Q�|�(������Z����n�=2ڵ����k�R�:��ۻ�L���;vw�}Α��N�߈����ٳ4��s8���'a�8�d}�@��2�5S�| -Ҵ7�j/p�qG��6TBզh�<��{�=�����ԟ�c�mHh�{ܔ�yӡ�Wp
�'��^ĥL��Q��~i��D��]��ޜ�-���y����(�z3��nP,!�Y��']�`�3�7�,�������%g9|�+������F� b��x�<��Xu*����Z'}pN��T�l*����H�B��$�Q�=�٢����ޭ��N�f�SW�ի|BUU�5���9oH �~U�J�Ύ���mRsᾃ�d�L�@��� �=B��u�Iyp�歄<}�T؁�h�%�w�ĲH����\����� }�Ԩ���T��"um;w��m�����&�7��Z��quS����U
��-�Br�%��Α�Ť�^T�SG�ÿ�i?�K��i����O߽��-�<�[5�;O8(/���F*iܷ����%�����H{��ؐ�������t�|����:��A��������W��Zi� @!!7��Bf&�mb��F�]ܹ�H��m�t�f���|L/��Me�\@�4�;�mCn e$��یڢ�diEۉ������.�W׳��N!��B���T��c>��fXpK�6TG5��X5�6�MZ)K�����,)sq�<��2�HPb�������������D��|J�������ꀟV�+�G�֋M�^/F�Zקئ����5f|��'U��K�e��z��ӭ��R��G�ЮM�qeP,���z�؜��/6�h��K�ŷ��D�Ft]83�)��a�� V���h�%�)ػ'n�w���CZ�B�؈b����0V�Ң���]�����=��G1V���6��g�_�C���֌Y�Uh�2e;3�mV��L0��p����KE5�e�3_�̄"�4�;�^�d����/+L�.�V��|�JAԌ�FJ��Ѣa �>CUu#�b[�`AF����.��ёw�C[��g�3�
�
�~!����&Cfŕ�H�pq�J}&~�p��hY$�&_��Of��s6b ����yd�	��H�����f|��?ԯ1���(�?~�.亅|A�B����]��,/�[�%��� |)զoI���"ct��T��_��ӫ���8w]o���X	���fIc�O�5㼢�U�U�)��z_6�߰��7�5���n�H�t��B��n�����Z,��S�լb���υ{Bu6`��8�72��^������wϨ�����8۷ʆ[0�h��]�,�kv��(�yDp�%��	,��=�M�H���CF8�f�\�I�rU�wvaw�5.Q��N%��K.�6��QQ�?u��2X��W�+!?GTG�Ǔ�ZJ��!��04�W%N�"t*���#���!�%��)�[6���q&V�R��{���ɪH�}	�!�F*�c�X�Gwi9�5T~�����߶mRT���1��J	� �K=V�m�oԣ��ϼ���1�p�Gf�����
�o$�oZ�hӈ˄�N��CV����X�=�P��X.z�����ɹ&cȆq<�nG����	p�(�p���NCT_.��L�ր�h;�$��)�ś�+
R@�h��u��a<v�`4�/WN�����#�K�)Ԅ�=ށ���λ��d�����@����D�
k)����G%ˏ�K���Ǽj�k��"��Ժ�>���̫@�1s�}J���:�@k��J�&+RAYw��P1�*�����W��-Nm������n�ڼ)�F֨��ݐsA��i�f���(\^5�� !22�aw���k~����f�M���ʹݥ#�O~n�k��Uʷ�R��d�(��uU��$��ņ�	�wA�_�k�;g�	��'N,�b��yE��%"���t3����<��d�4���dp{
$�5LI�7���༜�}44+R|����`��#�|yL��I��I���7.�8Y��V4
=�m׬Δ�!E�e/
C��2[2����%�$�d���e�üI�b�5�1���J�yo$Y0��������Ԧi<�QC�)�$���AK{Pg�"{6�!�~��8�2�t;g�.sπ2'��_Vht.we�j=K�p���q1����@�X;�������m�m���,�CO�x�������TM��Cbg�\�X������a����KV��ơB^i��z��<ua*r:�Tqڍ\Oo��o{h#�i"�Oo��YQ����?���+�������7�@�}�e.��=w}�����/% @�w���f-Q��~vyQT/>c��Wv�O�;I�ϼE�_
=���eH��Ǿ��1�(yy��L�"�l`@\��s	V�{�i��]Vν����X��66������]�z���Zr���͹�9�M���n��T4.�c�͌��W�l3�B���=j@��}�5�gr�v�W�u��ɮ�����{T k/�s�?��+�w��u6#qD��Pvn�`�|/�ݚ��IH�wnkҰ@��논%���>Um�\�@\8K�%B|X��F��=��ά��me�E�;��}��%;�����-V*?En@�rms�v���?��vNQ��@v� ڐ��,K�`N��-����{��7��-�#pK���b>s�C/_��7R���Y���IbL��/���'��a��yv.a�֛�!���������	~�
����!?&?"t�b .9=�nS����E�����c�˙�X
+h�^�j�
B�ZD���tT����6��M�S:�E�2-*Wȷs1�+ZsnR�$>}ٜY%8{.�[_a)y%����	ZC��A��^զ�k�%{tǇ#S�Ŭ�Ь���VT��އ�,/J�叓�J)��1�ِ�� H�lpW_c�/�A���7�=)a���Y�H/.��'�QG�8��}�5&o_���9si)~�q�R�{�v?�.�w���GJ?5�{�UAk��b5&P�H�]���Ց���V�X�i�P�}�y�n�b'�s#��������m��>B��u�.9��![W��D�|�-j!�>��<=�,7K� ~�UC�'"t{p��b�3
��ꮓu� D�l�P4�\������R��n�>f ű'.��	�#���W^t?�hH%�ؤp`�t/'z��0� ����@���B	�ͺ�u���@w���/-�W�_�����xZ��MCm�/ig��y����+��ձS����9i��!Im'�xϝ���|P�o��gf?p�am 7�C:X�
�נm�)]49����o{!��T�`g�uԃ��rfzL1�oĭ#d�'��m��Ў�	B�fv�X���K|��ۈt��z�� �٠�F�`@�%i���
x���S�����`�s��/��?�� �7P{���-����F ��_1sNj����o��vZE� ;��w�o�H�t�fX�Q>��P�-���K�|���.��� ́\�,��l��wh�%�̉�E������$`����
d[U�� /��);�2�jX0�ڭR��\Ϣ���WK3��fKe�Kv�2��Kck��\*�rs�+듚��Yً֕ͳ��[Mb]s����ˠ1B���E�Ä 5��s�����%G�Ey��hg��r��G��g�Bu^�O�.���2ɫpݧǁH�ًc�pr�s_����7\�Mt`܂���w{ωgU8E 'dY|o���TX?�E\��ư*YVӀ01�>]��ge[����M��%���H`�.j��909?����.���������BP�*,?xFTR��	m�X� E[�U8K�@�泖'�FN�=\�@D;�����3(�֌����)��1�w[*�S�~�78R�n�y�z	��h8%��ɐ�{��.���c�k�?��2�Fk��(& WXD/�O�jl��8/��P���&�e���Cq�'��� �x��L�H�)V���;6�|�%�qѩl3�-V��sS��R�9`�R��2������N{Vs���	J�}eEY�����R�
�!�7�	(���1�yQƊ��N��f,l���+�I��R	�=��e�V��(Z:#��}���z��n�p�5x�U{l7P�������mm靹���j�Z {�zM�eYҜ���Iլb��-�S�%<f��òP�𮃖�[���A��U�pn
`�76�ɘi���u7RNkn�R������su��Z���b������G,�����	>CG�u�j�e����n���ə�����ױ� �SX�K}�R� K�7��gI�t���¥R��7��A��xgǼ����<W;M4�%�2�)W,⩠���Y��,�.�7r֑mso!��w� @��JaC��6�OoH}r�!�4�#5����d�%ˈ��\j�����Z������vHV������3,nA�R�)��x �V�WB{�q���������9�5̽�^�>�ഡ����g�Q��0�q��Ǖ�W�k��F�@h���26��\k�do�z;�䗽�ޣ���tT�ٚ�W���L�eWk{�2��.u���V�؃�����t/�=�����j����ɺ7{��R�	�jM	%���}}U�����G��-�Za��Fy�H�X���@�';W�2���A!�K�sC�v�0�B�5�YW�s�w'$�#a��:91����Cm!0C�ٚ��� �nq�Y5o�#�0�jtT��JdW�����F�-�`�9=�9n��Pu�m�Yi�B-r����OL��-� ��l7OQ�K1���bE݊��y롟�k���'��Ai?����x7�,4�-�;�����c�ͷ���a�y�Bm��-9���B��$nj�v�<�d���m� _�B��o39������6��J������Z��ð�fB�!E��Wx>���h��)�k��8nq�G�Zy�{�ˑ���A�{���{�o��)2��)<B$�<k���(�2$f�i���}@*���b�5�&�@��XQܯ,I�͔ui8�啿�ߔv�Z3 �5.�����dM���,���}�������9�����v�����bd䁫�)������E�FP���GЉ��@k�m��F!}������<���a�1��ᷞ6W;��m�B4s��$�^N#'�Hu��x�@���l=.���d��b��W��V�b6k)Qt�}��;l[�ѽ���*L��A���/�+�\�L;�� ��:A�i���Q84�tOa%O(�fLSa��l0'ar�u��]���2\�d���]p<WQ�bd�M��U
�fR2$�`b�'�g�̓Tֈ^VTk���9��d�}�E��]��A��%���g��ͬ�b��-R�j����T�����̐��H���dm9
�BM��p<3-B��B�F���ݿ#���C�П�V��<Q�[�&xӄZ9�������fHQ���M�����ws�n��v�b�o�J�P5�sW�j0���U���I$�溔��.�����g5�A�P7���k�����l�������T���0_bqU����I/#�cB�� ��(q,$�!���L�/b�{
����I�
z^�ZpgX1��1d[	V&uQ�I0�p8�NmC�QɁ�) ��������잻=dK[����	����5R�]oU3��Xy�]��A�d�&0x��o*j��}IQ����I��)�@��W�k���uq��+LR�#J���~�f1��1"��4T9f  �+U+�Gi����q4�oє���ӿ��%9�s�ճ��$MW8�k!�lk�l���P����~n>����Ye匐yJ��������B�.�	"����c�.̻�[�K�<6@<M�@���t_��Jat$ܷpur�E�7�㻖ݠ�U��l�qcr����6	!���=�PQ�z� SL��K�#}<�Q��A׮����������l��>w9)}F�K��ǣ������f8�h����+�'"���U&!�'��	a�H��)�%�H��u9iLT�}֙�AO�Nv�-s�Զujs��ɖ��]�ɐ��iR�	z
��#�(nܤm�~������!�>)"n��{
 ��R�E��Yאe��_�@aW��%.}��ƶcR���n������8].p�84���C��-ay����3ƕa%�D��y��t�4,ϲ�Zͼ�a��0�g��R#�O�Mj$Zڐ�wTC�6�<xw����Цhi}I?U�u�<`��=fh=�����׻��#�������V�"�%�������z�&t�l�����,�q����;�IԇX���&�9��ʬH���U@��0�͋�u�
a�V<c��m# Z /W�jhv�*,�Ub��(E�J(�4��4?����C��)Ʊ�,�_F[�F�B]Nv�@+�����kU����ǆJ�������pģ@C��0�}ĭ^ם�B�,z�ӿ��\z��Q|�΅]�KO�~˿��&�(	�u��=�*6џ���qCg �d���~���mx����u��XͷQ�\4�W�a�f6���u\�O��v��y���e�`j��1�K�x�;fh��Q�Ҝ�$	�_]�uc��1��|@���U�ź����[Y"l�d�	�	��������f:��bʨ�eW6xz���Ĥ\�HO�!�o� ��*ts�TO]�}E�l��� ��y����j�ck���.�vv�(�|��+9�B������V�,P�ѵ���FNфV?3�/����ru�x𹂆LԡZ��Ә�xf[���Ԅ2��;X��5�6��a���fM8)���m[|i1ɲp'}�S��-�� 1�_�eڪo�wg|�3FM�����.ԛ�;��I��^���^B�?��5(�����ls���#,Z����ʿȴ���¤j\��ϧD�ڣ�� ^.�.+���
s�'�+��w�bF	vK��ɠW"�v쁉k�Y]��G3ڮ�90[�mg�[{5���J\;e��O��=2c�eU��U��_+�}�!wܝw��lӀܿ@E��
��Z�}����fՎ����anZ'��P3\���3X�/� �FK.�"�/���%u֞��V����>X	��yaa�s�P�Sq�����V$����4�?�g�	�U�#Q\�S��.�w����C��=ʇ7-�l$��M�&�шq��C���A�0<���̺��&�l����s���ڙ<jx��Ν��	���0X��ٓ?D/���>R:�N`����l]�2�^򎡏����,dQ��=�%��5�$�'����G��j�wP�&���F��)�YǯOT�E�i[�;n/f+�ţx�p����wSȇ������nf<X/�:�Բ��'��e�a�,��{��\�.�7����l����F ^(KDE���dujG�$�y����$�$�"׎z�����Dt��O�������1{?ɞ/|^��tZhq���t�����;Ba�H�f�+��>�aؚP�����?�6�s�*ݞ�w�5�W����4|80��OZ4o�����?闯�Q�ǫ^m��5�4��𬖿�H�Fݺ11��ݔ�O�`,��\<@���<�*,�}H���ʑN���$l�*|����(껇C#'3�t"���KL��Z����=�����-��.l�\��!-�8�ۮ�萣��TfE��*ju�8��4De�v����d�8
�o;#0t�a3��7�C��Rn�.�Q�a����J~8��';mr?H�	!IO����ЯQ�4²vq�+�+��d��w	��H�L�EE�u)���9�E��aȯ�N����gRz�
u�)tzd{����E�+&W�qU�(�H��n�KY��0��OF	"��d���>�����L+�����ϻrگԤ=���C��Cp����)C�囐��9���?]��Gam�,/���WO�?҄4�w{�1��{����S�Pٜ��#ZP���K�/f�xz3�FQA��_	���/�ũ8��K��^ַ�:-���"�G�ʃ��:����g�`�u5�W��{�V%�D躦��,��kZ�ͥY�rt�E��=^7���fcv��3K���x=5W��5)�_đ��ٲ��8(��w~�#�%��P.�j�G��s�V9P�@��4M�_>�k�ׁt�C�ƀ�$Y6R6z�u�_l��5a���|�Ԧ�C��5n	U굇*_h��ħ5&�oU�Fo����QiZ�40և�����ԅ/#k/�|�� ��5�@ɒx��@nN:>u��[�Ep�p%��SSK�X+>0����DzHkl�Uy�z�&k?/�2��u)'�߯s��/�E�>���w�pt�g�@%��摚�'&�j%?���h#����R��_�R^�-)N�(m�s���4HO_ވ?z�Y��ǚ�Wx�����H���~�/8�3�׸�ÅZ8VJ�S�3f���g->���'\E<-����*Z��	)�YãH���ib���ol�9FX>�^Ò3��_s��Xѯ��'�k�o�Ȉ�2��$?e�)G�����'C��Κ ��8/[������A]�2�a��ro�}	�\��7�m���2�>]+�Дl���̽�=�б=H�lh�M��-h!dΕ���4;C��Rjn��%���*(�ױ���l�ڑ!ջC��JR��~�O��wxy!-��6�<�f�\�XO.w��� 9bg�qy%��aK�(�gaW�q^:��p�#,$��t$C6�#�>e���Sll+�9B��C��hI�2�B�+
�]�zj
Y~*�ߠh.���Ǹ�����Ɏm���)��.����5�6��۶��s;l�
t��Z_�w�P�F�@��;<$_�x�2tG��r�bu�v�$��ҜM2�-ia�5��
�h��j�9��c����c�㡦��_P�ޙ.�ǝ���Y��ߓ��*/;f��`u)y�i��	]�Y.�3/�k���7����"n���l��I� z�ٟ83�]8g`�Z�*�-B���:�nR������u��U���t8*�#1:���g}+k�肅��eJq�i�`��]��G8#zX4RHљз��%�����4��?���6;�Sh�PdÈ:�7#gW����U�v>��P��hy	�	�k��A��*l3�q�8
�v���a���9jnҡ%e
��2<��h3'|��үN�3h-��K�G&pZ
�Oĺ!3���}��}f��E� 6�[a�d���~���Atv'Hh{��M�#՜Ռ/|�HZ-�
�� �4�H�v�� �C���u��QS��f�b�%�g�44��;��o �Y��B�����0!r�U�c��Z�n|58�2� ��G��<���f BS����Jիq��SQ��D��P/��f'2v)��}���gl�0c^s]����EqIZ/.ɹQ�kJS������������s�-�\L^Bڊ�8�X�h	�}��SD�Z{;��!jf��ot\J�
ӯ�^�Fs�zf,��­���GA�l��-G�  ��&�t}l�Ba�c�$:�W[�h0<���fkd8Y����n�@7���ah p;X[��y�ې-ă_3�""j�pE��ҙ@���_��Gp+\�*-�A0݇�{��|���G�_�=K��m{ZK�,-�3��:��'����=�,0�xo���c�CH�g
h����X<�f���`�Z��O1:C��*�%�o��By�a�1�!R��IP�1iS|}[w%v��^����y�yP]s���㭜<䴴.���>�lh��I�нd_y�z�Dbb�3yʓeS��k��p��=�}�/��rA�|�ܝbP4{�I�]L����Ϊᦞ�$(��7�W{��\k䤱3Xj �ۆ�����NM�&����K9��[�÷#��ׇ������e���\�8�����9���o�L�tm"��us������M���gW�A�)��b�<�0d:�D��SZ�,R��K,����U���E�d_\�(��+�Q�	�aV��R�:���ǥ ��o3:ި��?!p�����RUc��(m��ph��7�R�u�
��K�	ƉU@?C%��� ��X��S�Ԣoհ^Vii@x�M�k�dmxԝ3h����ZrhUy0U[M9��l��Xn�s#����c�UɈ��K�F_@n�IYj)�-��X�k�V�;��kݚ���������3��.j�3��L���1M�ۭ�KI6x���65�ޥ��ne�8���K�s�0�n����ma����<��':Ů]�:ܡ?�m�+-����@Z-8�k+�8���_؉��ɵ3ӭd��H��Ś�hb~��N�Z+:��G,�J�g� ��(�'��Sh��98�eCH�[y�s��ANK0I)���J�.��Uj�N�t-k���@��wؽg#��@�te��F��|8�'���Z���Vs6����(+GobrW�T�R���N�JL�Ӱ��n��Ǎ���`����6�ZF���Kٕn�"�r@�r~�X+���o���5�}5��^�ς�|m�J��\n�Ǥ1��S�fv�h'ӏe�81������)���am����UҙF^�'���ǒ��[��0�6>�)�R
V3��O�����+���F������O�FCy���Y!�h���u{��`܏����j��.`�n��,��q�h��ˢ���,��k5���j/��}&v���#��h
��N��_������(q��I�<Y�W�}�)n�Tf�k'>E�p��S?������=3?��fC�c��dG���ͣ���tI��̉Ή��}���N�B�O� �:�f5�W=�3<z�Z����4�ڹ�ؖVT�Ǔ	+���BI��}�� �\}�M')�l�:<������I���/���o�2(,�,�z��הp�nF[)`A�FUu�ר�l:��R�� eʇ�9�9/t)~�4�-��xPf>�/o�Vf����n���[��,���ǪD�g&Ic��A�Qp�k�)	=>��8�H��AZOT�8^�dj�a�ܘ��IJ˗a�����: �a���j,�ɏP!(��^p������0(��Pc����)�������"Yx�L�%R(�\W%�m�� p�|j'W�u�U��sG�OD_�ӻ0�Y����j�����5NԜ��7qǰn�b���Ƒ�0�5@�V��@,*vQj-��%
TyIW������^�Uwx�WZ	�� ?K�uҚ,����+SCcC���/LI� �]�A/J�5�9�z8Y5�%�-Z]߲�7��o��,������i�����B3֡��It�p⩠�jj��`Z�?�L%Yc��ؒ ������Z=x�Ñx��zw���»K�oԤ���O�o�i�,\�?Ӊ_y�*%{����ͽb�
�%����&b �־�q~�#�	:-Q�fSŒmC(,��:Ǹ��[�C����2��DZ��O������B�/�K_�/09���])�9>�T�
�ch��~�R���96=�N�L?WS��u������떤~TԮ+���T�)�D�S)�'���o��Y�!R���E��Bŀόryw&l��8P��u۲���j�DD�?�
Dՠ{��%t8��S���ݸ_j$^���
n���zP�"h%���K�ᒮ9�$ ����/�P��x������e�}�D<K.ل)F6����%�\D�k��w	�	�ۘ���J��V�h�k��˒ �Վ'���r(�!�,�����1Ѝa��0D�����<���3�p�m���'?@zD,�G4=��y)���8P�H��k���WT���&��-��/�I���V��RܛJ���������<e���΂y�K��.[���sRs�E���$p�(�/.�䄶�l�a�IRwFq���H��4H��Dh\�$ܭ��NO��:bq�c �@dI�n�}Wt�hZ�\�c���y�bk��N��@%�C)U���O����q��T�A3�F�h�'�"JX&~���E��d�W�xu��np.�E�*��%|}M&�Z:�NE�u�t-ʻCL��rg~t<с7�{3�i�T�����9AݸW�]��J2)~F��yⓀ��`� Sf�"���G�:��j}u~.��D3d�$O#�뢲�2�<8���y3L:��.��̛@��F�$:��<�����T�qnФ�7n�҅�{M0���Tv����o�
i_X���2�?�n"�:^vxVd�*y�h���nAicS���%X6����>�m����:�|y������L�U_%������e���L�5s��S��5�O�A�9��qQ����U.��^��_:�&[N���9�	<t�kY]�SF!��MqE�Np���y�RP"`�3�o�")�s����AP�3M�s�}�ٗ�:�ԏ?@n��=���Yz�3x�z����R�����l�k���h����W�]�`A��)�8|����c�[4���^��������Eb�����VN�g'[c��k����M�<�D������#�\�I}���ޤ�Ďv�t_�]���zF�%Qp�8p邦l�0�R'8�I�`��o�ԋ����̸\ڕ�c�ɏ�C�u���Y)@��/h���d�jY��_�FeI��N���c�6�Z1�qC6F�]eL�f��SĆ1�W4+퐮H!:��.����5�����!}�8�]J�x,^C`;�J������7�D�R�U<��͡*@D���ے	Y5��b v����^PLX��,��vCp��\���f�>�ǘF�|b����oo>B�ΜW_�5��ҍ9�d�4!`�u`�r���v�ш#V��re?;R�j�T���$�ܺ���!�C��$]~u�2���pB��
��3�X�2��g,6H����G.�_���'ޛ��|��	�+!��f�!o�fD� t�fbռz���EW�<�PY��N�E?����-��W$Y`*/V@�hy�u�{�1�x'�����aN3�f��
e�0��PκԺ� ��M/�g�[�� ���i��/M;G��I���D䨕ӑ��y-�v^)�M�&�+���g�6g��yD+�H�B\���<�F������M3[���a
�6h�N󌀉D���迲H_�=��̯�h�W&�Y�"pq;o�T��q��ۢ�٤g��(f��B`�xi0�M�<����V����[BN�|v,o�nZ2�P�`i#�ås�D��x4�'��I�k{����t��B)	n���J/���K�iͯDI�k��l�4�H�T3�
m�B�q�d6ĜT;�qUT �~�٫Q�F�x7��+{��#,42k2]�u�-�޶��>1]����O� �����;�E�B����Br�wO��1�~a��A�v�ۨK�Q�]�.};#F���
'�E��F��쨂�Z�:��Äjw����J� ��SM����f��I�ţ�
�PW�UP�řD<!���~:WO�Ѓ�C�tŰE�ƚ�,5�S�N�=O�f&6}J�r��L��	��'C�γ�^�Ф�)3�~��CI��زY��r��m�ZVQYY"���9�����b�T\ 3������}."w����e���Qx�,2>���Ae��������D�癃n݊�Q�;N��RZ��ʹ��h�۪�t�Ͷ��Υ��vP��њ<��gHm�J�{{�J���n�%��"A�'M�q]���N�=�;J����h��d���:�G�Y��Ŕ�i�y��bR^�^QkW (�D�]�M-{�p-Ѣ�Ҧ:CN�O�uŹ�tJ���M/%�S���0)��KwAt�;PJM�����yF�Q#ᢑ�c��>	���ʹ�Uv��줈A�Y��i	�s�ptll{e��e�ut��5kS���/�� �HV�Wn�~U��G�-��!+�`�����m�V�ݼm̍ l� rnɖ�T��w�y�ĺ�j��,.SR��v�.�3e�˟TLk����T�2R��9�I��E����JX�͢)�r2��e��_$���t��_n/�i�Y��s��˺�y�;|��A�w�"ܲ�����52�W�L^U�a��	G�Y���,�����
��a�O`ј��)&�]ψ�)(�`SɃ\ڜ�p��V��Eu����#Sl�Q#@s՘��:^Z��6�<4d�j,h[��m�f�:u$`H���zv��on�a���E�l�{3旷��K��}MLǐ�_���4M�z��n)@��(��,ac'Ҩ�%�� �ý�^��}$�fb�֭����z�E������zQ��9�1�c���J��q�+������Η!��:�C�5c������Vّ�ퟝo�T�
wN<
�q:(�0�6�|�1>ɒ�w�ө��������YjZ�-o6e� �G��2��J�~L�o�~M�pn��Q`FJ��b�F�>m��EC�!�ٵ�<�R(�:.y�O���@�-��|�]LT���c�s*ݻ�����4�q��T8w����>5�j������BF	���ͨ�����9����K��|%�!�!p��-�	J�����`����C����P��Z_P!�B���
�J��H�I^b�s*�
Y����vG��8H� "'�-��V�&EZ'��FR�YV4`8,A�����^��7�܆ʿ�w�+�r�X]�<)���2�z��4�㌩��>l�ClC�nKO��OT���#� 	��ʫ��ޑ+vjlV�v����rT����.e�����Ƽ) �ҭ�d[M{�u��x�g�����g�h��1o
zq�jh��씠	����?r*�O���j��lsZ�U�z]YM�k�����o&3d��@��+����ZN��V=���CBH̉�g��^ZZc�5+,�A'�۹iʵ��>0'p*~����5�;����>�ڊ���ve����,��-�j!y5��|�UCqd{@�S�9��U+I{9"��^)u=!�5w��[ͺ���?S~����|<}b?+ɶdo�	�oԮ�AYL�7�r�}��aO����NYaO��T#O��^��1�sGOP�Q~��!�av�S&�~�M��H����+����p�������se�G������I�A�Kxdj����n�_�?!�Q�ꂩ�Y���[�[�Ӑ��u_(G�IV~��{��śc�J�táװ+)Z�;Ɯ��~�����s�Ϯ |I���^�`�Rc��5�ʘL�z�x%����ĲNI�O��l�Zb�M���~sx,��D��Py譤���._xD.�����|��ǌ��ѭ�<�S� W�޹#�2��"ޭ'-���jd�Ĳ^�������y�R�6�<_5a�6z⧵�E3���Q'�&v�j����aaL�{�.�'����Z4%8Q.���.���Q���@���a]���I���.Nҕڶ��n�5a�fc\5 C��A�Iڥ�31�A�y�ȩpF�C�G�� c���Ď�}��|�Pj�x͔�l\��O������cS�w���Uw.�z24's�Poxű�����G�f~�@�u'Tg��g�}��,t�����Hiw�gv���[�	=H"3����[�\�/7��X}�V��I�n��a���x%�7B<Ay�8殌�d~���'����Xv�S�R��<%�]�L���ٹp
�ȶf=3)��1�ŊI�r����0'�w5 �C���И�o\��<2����R˔��ߌn�9�)��S�G��\gj�t��>H��oS�@�ܴW(#;_���]���b^^�r$(Jp�7�!�� LH9�'摄�7�b#2�E�-l�\�Cv%��{�����h�h�U��Z%��t�j ��@2�;���K��*-�Qh�|��u� :�S��+����$ɼ����fA/6q����=�ܽq�ۊ��&��^���/n)<E���b.����.���wǗkR6~����:��(Q��G{��'m���@�@%�[�=2	bR���~����-1�M�i���P���^��8eQd�֯�Kɥ�).܍!�U�P�~.	���Y�8N��Xvc�Ė�9P�(�n<�^L4�:�;ϪxɮR�5�t�%��ܠ����������&�L|�1M.Т��k'��V�޵eLۊ��[b.�e �Y��5�1����
�ps�}Q�Y�
���k�l$O�{��c`f=�s�`�(hϻܰ�����06��������PMx�˝+��a���P�����y+�]"��5��[ݾe0�g�6��~�-���R��
e &t�1^8���j��eI�Ȅ���4���owΗ�`ˏpp�F-,��� �+l��-|𐬥Y2�Fx�� �ޓ p�No��cg�]�t �3r9Y3�eJ_U��I���MG�����9�dp��@3Sxm�IIٹ^fq�p
-�].l������%*x8�=�~����Z{s0��Q��{ь^鹚�F�%(>ݘ,�+K2��p�ƹ<PUo�MR,���]#�q��OY���J8�~ɻ׽c>A~��	���Unl6!H)�$7ua/3-!d+-���>)9"GZa����ѿ
G�A�͎)2��cƌ�Gxu�`�h�h��cl�������N���tOf���G�ɭ��ЮZ�qg����9I�[k;L��v|�J=2ۀ���6��+�A)$!�dEԟy��HK�)Pr�L��cuf��2�F)�W@*�CƎ�'��$2��������$��S��?�ì<�b�$��L
Fw��>ȕ�,h�Bie���y��!�AA���2��-bO`ϟ��w�t9X�ζuT��)S��ꭐ� �B��� �7���\#�8Ʋm:�_-\C��k��I�A�vЋ#����m�APњ�"$���k�4��4L��]sq�i�cw���(�a�����淰����?]B�����o��T6��y�v���/����H��7�ӷst9�AV�k�;�d�p�3� ���&��|��|JF]��¿zb��B[��x���X��ͅ�oT�wܭ����wS�b�!���g����`�`
�ȷ0b"9pG�/�\��0J�Y��_��৶��rXHfo�FY��X�o��>ن/&���� !p#��䰁]�0�����$��N�u}Q6�Ħ��|�u6�A��g���,"����f�>~��;����$�e�0@��˻uD7��u]kA.*7��s�r��-n��y{E�~�`���	��P�E���lgM�2ѓ��2�2�r��=2E�%�GƎ5GC��2���'z��=��g�B+ -q^�A����y(&E���T����f[��$'x��kd�8J�x2�2G뢁MT��f�)ׅ?k���Ԡ� ʂ�\��bu���19ܽ���~ R�p�1�����ѽ:$���j��Z�a*�ʽL�����v�U��D�$rƲ���M�5/ZH�@U0<����Ӹ ���}w��w��5�,:o?^�^i͹����4�H�4"W���F2^5)?ߌNp�����ۋ�)�qk����%Z�ް���=��^�c����
��J�")>?�[�#Z�{�j�O+���]>�(���N��N.�ګ�z��\�w�Y�j�P���ٌ�_��=�(3�
�SW8��TM��r��v����"!�`��ΊV=�ស��e&�>.���������X+C"E�=+k��ܢV��CX�/%��Y�K��Ad��No< �V�(�	|@$mi Ő�̋���?��6���N��Ӳ����b(�2��Rb�+g��t�`�=�	�I1�V��*f\��c?�T��#F��8�����<�0����{ⳙ�>�j��� ~p�<���/��͹�$bIҺic�*�=DV�D���n�eB44U��>�����N[�]��'h��*'x|����@	��&wq��X�u��.��!���D�W	��p��*��f�A��P� ����:O��r
V�a6|â]� R��f�%gg���;0�'�P��;S+=#
o��ez��*�xc+�OB����'7w���������$�]�(z�d-u���42  ���["}�<�!3I?���36�n��љr4�M����^-�S���d��;������3r��U��R��S|}/���\^����zaѭk*��w�`�2*�����2F��XG���kOg$����8Mt2�!��?Ç�9��X�0�!W*q&uuW���_�L�[(=�\|hl�Q�[}�����碷�d�=�ٶ�0E�3,����Q͚K����r̗-�{�i_�Y��%$8\���c���f�M�P)-��A�j�il��[�����s���o�1����i[v<e�$��i��9�������OK����n�Շ�0��R��y-*���Ȟ �䒔�� ��I�ik~l9/\�����}*��)�˓�=�T{Ղ�=&Q��ћ�2$@�;� �FumB��P��3�:'F�r��f���B���������ZP�uL��C/�Ф+��)+����9�c�*��D�lv|��Ň��gw(^�M<i�7��4�Y1����󤂊���D�'ɶ��E�y+�UJ��1F��]$%�Ӏ& �^��^�R��/zM֝�QM�Xֶ0W�S_a���g���!��]��1Qq/2h��b�K��Hq�y>�O�H#&ݡ���"[�J��z�Hb�[�"F&{��'�#u���TZ����x˔ݮ ��wL����W1�F$�Hz�(���/�;qQ99O*�U��Q%7�(sW��0� y�zv�����J5��8_�QdU�L�cJ�_��Wk��r�����-����c5F�
�f��D�?*����bq�y�Mp��P�J�;f�g��eYH�-������F�pdL�g��G�x����K�׹�lI��,��h���60����I1s��N���`}����6<֤C�F�|T�$�B��P�T-��c�6ڱ������o�=���.����~���PO����°2\��i}��������B[���CX(#������|%�,����C�6GOź��sE� ���L���">�{��+�p�&�~�S��f��M<��Ȁ����K��<_j~I���1��sǱK�ңP��0��al�b�;�<�='�� e^�G�l�d7�i�dD���������T= ���E�1%��T��(�nX�7�~�/pWg���o���ܧ{����D�ȭ���S�>-:�n	�"\�!Q<q�)����_�hF��7����2_����)}��˘�=/��wp��^�pp��ԕG��!�1XH<��	=�I1Ň�G
��g����l_�X���O֚�/���h�ƞhhuyw��%��%1܌S�	G���{�<�K,��Ki���AO8j��`2
����[5�o&�C��vCL�|}�g�nLڵ�+_�3O�]��e����uG)_� &����qv)�wU�M'q/��9��^���Sb:��1(W��������_���(y�\���iI?��<��(�{?`^o��R�&(1������)��T�;u��@k�=�NߦR�l��W�b�u����ЭD_[��yi��붯k4�Ӝ��Κ��\-M�H�<�"t���"��57�*f���\��pN��(���l�!��̯5E�}[�5�`P2s�h&��}��f^x�T�����v�!J�"����r�;�ZͰ���I��*(����?��U�v$�Vѻ��Z��R.�9�ձ�y�����Qz��`��?��ƛS���Y/v�[�g�z" ��a?�*�:}m�.��[�-���|������kPk����7-V�DC��ڵ��ē��Sd]f�=��	����dD�kǉ4��>�ʣ���Q̮{p����t$ׇ�q��qzy�����_�ߖڌ^űi�g�ާ�Š*���G�v���>ą��Fu7�JW#a�P�߃NŘ��5\e�'�k9�B��F~��=�T�D5���l<˴��wxW�&3R=��dŲ����<��ǃ%k��Ʈ1F���[??���YwG8�7a�I]j�Ӽ�I��[?���L���rhw�S�s1��f����{�T׿�rF��34`�<�H_jՑq��n�J��~�4+u˛�%����C���u�@��Ax��N��)��ޤ����C��z:�ژ�EC�:x����,Q�;~w����<�a;A.���W�±����jtPF9�1`��R9���/l�]��@F|Z�y��(�g"���W�t-tN��(s	�)�n[����C�n�r#ٺAͣ�>���K����@֌3Z{�QzŖ�t7s�n�9�_'��VC5p_��B8���!�<�����m>C��-?E�]!̿R�����>���"
f�RPzikz՟'����%4�K��o>��.�Dpz�N�D���J���WB��|�5xPh���qZ�;�7��}�����,��.�Z�P��F�ң&/bt��&�o��{	fO=#%�����yf�� J:�������H����K�p�ytjB���ظ��釿�}�x�A�C�o�jj�"�ց���&�aqݮډp"ϓ�m��Ў���k؟��D�� ���X,d�1��SМ��9J�J<��:<PT�Ȍ\�7aљh|Rg��W������d�f+V���*ԙ9�q�(�P�*�4~�_lu��R��Ǳ�K�`l��t'	h�B�F�����$Ӫ7�6c�p�E>2�T ��
���]D��tc�i��f2A+��i q닞�xH���b�]2u��D~W(X�R�Q�2������m����K_u�C�|d~:J�db�ob���C��6�ү�=��jt@�#}>�+3>y%�1F�)�,rn)8���2��py~7]r͋�9�T�t�r=4G,��\컁^��>�ʙ�]m荫��h���MYE��NU�fθE�J]��kc$�AW�¸m7w��$;Z��Me]lx�@mE�q&�/n~NVԾ�5���Ño	���Ʊ?G	�  ���m]���N����;e_$p�G<z��p�������i�F�Z��v%�Ƅ�<� d|����֖k!9J����H���5��� 3�Dҧ|1�u����
���S���4������7K����	+0@ �S!f�q���֫��>�qqk�b��:�ﻞ>({�I�Z��e�P��H�gf�%�0����`�� ����U�}�#t�΄F���*������nħ�-���i�������}4-���z�J>�ޔ���.�rSHj�w�<�5$NB���N�#s��pd�;�y�Ż�(o(H~E���

`�x(Z���(����@�L�ɤR��U���@��^x<@a���V����6rb0,z=�&U� ���.h.�i�0���Eq�]�}�a���rC}� ��Kr�&U�ݹ�F���c���T^kv��v�ǥ�=���yV-�2`*]]�Ӛ4Z����.bp1P��q� ����4xi���&���������3��"�<��f?��ES�(��%�m��@G��-�[��F���A�l ,0�X�
���'�Gy\��_�mպ�,���Nw� H9�ҹ0�S\�ֶ閄|�˄D_���}��w�����@�4���RDO��k���1V#v��I��,�����V�P��F#CZ{߮�I{{��5M��_5V�?ߦ�?�'��yqc���9�Qd�����w;��l7���e���L��J�,�tgt�5�Nq �?�G��t�Sg��!Z0�1d3�<a��V�F�ԧ�Q� e�� ��k�U��J��&��2/O�t��|�̀w�\�'�e��ݑ($)���Zo��r����NK���<�C��]�mf���t�萹�&G4N�.ڿ����Gd{q�'P��w	�ir@q.����T|����Y�v�ftZ�Wx���Pj;���<�D�]�����ۛ.�r���[�����{���(�~]8w�Nq�s؞ao!��,��CM��6���z5�j��Ol��W����TF�ݘ�u�f:�ǓK�YyD:���dy���}����sF��V���@r��|b<���!���# �]���>����TV������Cn��fD��5��?�zߞU��ƱS���躡�%^ށ��0�/{�ۛz�U���H����X��&n�a<9 _.����5���Ԛ�emtCW�#=����ϯ���[O���)��y:JW_�Uҧ�&?�!�!T]��eg�R��Qx܃cS����i�lFBʿ5��Fɩ��-�r��(r��|ȍ�ր�c��I�n@�)���XW�"`�s󼟢��y.�ȥ����O�����I�#W��±p�{�%�����&�dgt/wr�W��x� j�������p��{�T@
�-b�P*`1�����jr��a^ Q(���D�L7�'�wdEk�Б����[��U�ijވ�t�80��[���j ��j�~+�5����)���|�_��GJY���V�Vp�_BL?�=�����SOg�2�W5p殜��4�Q88���?��{�x�̪�$8Ǵ��s��o#���|q(�hۢ���]�c �o�5q9P�K}��}���5��@%��$�Qq��~\_��,p�=������`�νҵ��HN���IU�Z�5w��Pٸ>w^�����=0���Wp���"�܅��|��dS�i�:Sю���N��6�VU�6C����X5�+M����)��c4�����X9�q�ZQh�#(�R�H-���x	�-��1G��K�إ�ݮ0�V�A�
��u���m��@��q����3�O��<��	��\V��}y�cm��ՉD��ck��J���s�2�����M)"E�Y�XAE�EL����Ҁ��<3X���=���t��8ܰ!�I���|�������.�dIO].6��iO�� �D}$�1DI���=G�u�����p�f��i��c4/D�1�MczeG���Qͯw.�B����g!g��֝d͐��s!<�%=�vċ��@c� +X�x͙��8�^(��1�F��tV�w��P����|Rv9��̚)'��=CmpQ�EW��r��i�����|����o�k�C-3��uro��i���H���i���j%S���W��������&PqՕ"��	���$\�z>���X��e^c�	§@��IIf]B ����N�m[�b�y0\��%���[�0����T7~/��~���������~���������v�'�")@��F�<�%ۃ@�Ty�,�X��&J�Iw���7�h%�[y��E���A�ב��^��I":�Y�����y�[�i4'a�x�C&����߸�?c���h�q�&rl����/�+Y{
��h��ϣ���J~9 vE�*��&���B��R}���8B�:DB �Ht֑���&�7B��\�0�����v2��&��Y���&�����y�O��7��i�g{!ڸ�<��3w��k��oE��ތm��t0�G��s�R'}^�x��P�!v�t�!��9+]�N��
D��
�N7,��?��NC17�
�[;��x�L��A�D�36v߾E({�>g��6�� �c�}0�솞�����������N"ƛhC'�a�hΎ�yC�T�^�UP;��k�>�\���:� =F}�ސ�y`+�h*n4}��b�/y��Lƚu|�p��H�lB���_���Q��B�����C���~WL��!�o�.pC"�b�LD4p{*��;=8 �I�%uJ�L>�b���S� G�qm桴<�Rp����9�����2�1���-��3��	;'���j����u��o��|�W�b\k�lӅj~��?����e�YBE.nrj(jw��w��/�����͆5�zb�=wH��Ra�>�I�P��&�o�*��>�2_� �tԝ� �Y豰C.:�ͦ��o�d��H��l��Z�Vfm�G���"ۣ.Oi$4��� �˚63����%��%Ul5e��פ߶��HR��}L��9$��ڵ�~7*����-�-�rٵ���x���.�V3dEcW������ԥ�S��I�O�� <��sDۚ�ɟ ��fEK��RF�O���G��o������.&-X-�p����U�WZGc\[@�~p�wx��U�s2�sfRp�,[�v�HHO�=3�K�K Q��k���n��# :>��F)�2]��:�&kڜ���wweRx�4K������ܰ6ݲ��B�|h�n �\r�$t�N �Qi:z:)�[RIi����O@m�-*y�dDG��i���YD�2�� ��Ei��Vv�\."�(�U�l=rW��2Pp�O�:����t�<[�{(�|[ú~�繤���f6��X�w%�����oWJ
&���O���豉�ucx��O�2Ul����7���w�x�*\-�u�DG����nu�h`�ݔ�r�!���2g�P,���}�Ə��(�����c9��BP����R��!��}RF,��,�1ix��Z�`Fnr~t'������{nW%:��;F��rL��d�+�@���0�Z�R�hªf7N�۽k���c��P3J\{Ԯ���=g⏤�,���^�Zhr���;Qd����	O1�|l1f�H��
�u�-�
�� �[ϰ�|�hw$c�� ����n���3�UMr�Ɏ"��yxA�x�φ������w�F�oKP�M�	M7�'����O�`���,ݴ�k��HeBL�,�M%2���2�ԗ���SS{P�ci���5��1��i���Gί�"�@n0�h���R ��Ky���b�XEq	T�pD���.�=���Е�E�Kk��j�DCz�=��C��9��HFį{�����d��T(>l}X2g�񃬐��|����G!h&�3����vkf�u�	2��4�/0�8*d�j�	b.��V|̀7�N���ƇM.��6յ�=#(�I<LjǠC��gq�33i������ġ������;P�f����;/�}^���$��G�����]ѬM�L)�ՙ1�������gD��D=�QRpa���R ������؁���L���r�����mY=�&ǵȬ?Tl ��t�6-�|�3��_״h�(��]:��Y�(}mk��W5d��\�Qz0%��Ϥ�rA}�4Հ����zo��=4)'��n0# �i��\�B!���+Ol�"pZ�^]��a�8[Q��Yc9h
>?��,�z�K���'�j�mA���V�����ߢ�	4O���Si�����f�pX�Z?Rh�=� ��h9䑞bc��'��Bqi�(6�Q�I��:�=� Jp~
{�o�V�S��EO�"��X]OO�h��2�v���9qE�s�b�+��ܡ���h$6z���6��u��Y@�jgzs�j��[���"��	,�{rhx�ds.�~�R׎�sO�z����,��;ik��Ş6���I ���γPf�P��	�`�h֑>{k�5�p4e"A��B2w��:�����<��=�z�D���6 ��0��D�HfW�-�[�P��e���ui�H���2�&��S{�Ң�8+��w\i!�\ںb�DKߢguZ��t&�eZQb�#�,
Z%�F������SO�P:��d�Y�NT��ԅp�����@�}�8Ns?%�gqW�z�^LG���0z�WWl8�;r|��&�Ko��X�o�J��<\��k��Vy�u~�z��A����9��c�����MÚ\h���/�;�Cr�=[}�,�U����3�1i����Ĩ�v�6ҳ4j6fq��a������%�.I�S~y���u�#��u�[���Q˖A����ƺ��(���0�]��p�<��ƾ�c7눲��N/�Jۀ�y8M:OCty�~þ��^i!#��VV]�FVv�z<��,ҮמQ\6��>��H*G���/��@����M���ȭ�`+m���)K��j�R״h7��IT��n���U��w��:����gKe[��J	8;���s6�B�?GJiK�(���L����]�����۩@l�<�/7=Mr��(�G�F����2]�#���5�O�Kڕh�����·lYO��MmQ��o� ����]ԡ��e�◵�;T�b5��!O�g(LɛT5qۄ��_��Nz��e���� ���E	rb���
�A�K��*hPj�l(��^!	?f@N���<i�ڰBz�-G��0�ݾ3NY�;������8[�=��$��KDT0�^/�MW�UՂ7�_.'BzY\{��.��������U.Fu\�\���ى;q _*|r��2�i�å��$�9jl��ލ���%�6H�FDu>�1u���-�[jPڐ�V<��q��;j��%Uy�ꏿV/>>�.��܋u�z^��OU@�/�F���tZ!=֞�)㗼�K�b!Y���V0!�X������{�5|?M[�A0+���>^r��!��ǯ����6� Q��=!�{��	h���TPx�6J��:��.j���y��%�ލ/Zƪ��7��©@'���CO�-Uu�~��
ҍ�j�o�n� �Ui��K9���L/�COJ.wp�y�n�c��x��e@~5��'��[�����@ew3�d�2^W-&	�RR�����9~��yv��/jQJt�4o����2׻������!i����yA%pr��m�y�WR�T���:��	�C���>���[��Q��0i�{�����T���*j��W��U1�AD~Æ��.�'Q�P���~Ӣi��_1��q����@9p�[�5!��#�Q��Q��$~s��ܑ�Ȃ��'<�O|r(<ܬ	����K�߃$Q���W~L��NQM��4;�HL? �Ȕ��Q:\�%���Ũ��"��]&�#?��'Pu���j��ש,��=�����TS�qѥxװ�H$X|����й�{N��M�o�n���8����8�L��7�Ҁw��(l+�<��R��w�!�t=-=���hG-����c\db%>n-��Ca���[�|oI�Ht"	F�;���������B���7j9u?��S�9i^!nCy��
Q��b�ļu�e�R�e�է�g_Ǒ6Cf
&�{W���>�N�WУ�?�F$zXXĸ�H���y#���H�9�n!��B�NbJ5.5t�H�u?�U�Y�QAF���Y���ݧ~����)�(4���P�!�b���ƻ]Zx�Q֙��<m栂"�$(�y/�=R�#�ܴ�_�$c���_xG�b�1�\�B��}��LXm1}��^e�^=9�οS�0�������!�9��4lqDXY5�Ґ�M���_��}D2��*��\��"��͟'~�>���~��h��UU��kZ��g�ѝDO�F�rp�<����\�������2��+���NE$-
s������WV�h��{��֥��,�X��ƛ�����0M�U|�?^�E&L������\��ի+�������������L�l��q�iD��;�{;:س���\}㦭ҵ�Xe����S����"_]�%�]�,�ta;�K���M+A�!�a��(v��MN8r����vҬ*p���G��Fl�z|P���0,ƬC��/���?�U�l�˯f��K�!��__� �>�(&H&B6P�xɻTRg.7IHϮ�� ��W�M�B���� e�yUrl�p�4�[�H*�'�Y+�� #n+��(�I������7�v4(������o	䘮O���N�0Lg�{�f?��6�n�(��I�1�>O���-S��;�`	�2��׆�E�5DJ�b���ƿ�B�׏nк翃�<����mB��7� �><�3z	���4"�D�!X�� ����Ȓ���i��}��#��e�`fjlj����G�  9�&79�/+���?C�+*̟HH�.ļ�q��T� "_wS���ɕ�mf�ʡ�|���q�q��rԷ7���2zO����E�=)|�]h�q�����J�$������s�8�NͦP�9�������.��V�bB������k)����O�)��ҍZo�0�������<�JBmh�腅����3W���v,�m��bK;��I�O��Ϛ[E�@'����A����,E���$�z>gq��ήeណ�_�q������w �I�|�GwAr6�αUa�?1G�_���g �+N��5	+ϡ�`�_��Ӡ�V�A����n��!"�u$�޳���J�{ʩ��M�y*��'.��G�&��o4�������Q�m��Xp�D���W$�_f�}/��s>�]��W����O;O���^���1w3���l�$1�zX	t?
�#��>���Uh��Ew�����+�v�9�=��9f�ʲ� �sڵ���Ȉ,Â�'�a��oH��f�>���H��)3nBw�J��L%0SE>���$������{�E\�M��4��&:���0).��n��N��{���ѶfrG �+C�o�^,�����M`�n�Na���|q�Ou�t��[�!�r����I�B:_N`g��ːk.pU ���jml	�c]��h��F-�*�I0Z��5���h�oo�U8���3M#�>�{���"���r/BS��\}�����]�$�"a>ڎanH@LQ�Y��J�ҫ�tR6��3���Ƴ��A�-�Kț�}��oۇ)7A��8�?�y{MR8�t�5���)ZﶰC�f���7����J�S����q+n�QAY����w�};-�ۋ�Rr��H|�����/X�0�2H~~ȋ�_ 	�W�ZXp��퍎f�;�9[��A	��0���ꖇ
����U<���d�GږZ�����Ы�V�Σ{������YJ��`1��3".5H�-j��s��wݕ}�X��.g~�-T�I-��] ��c4�7��a�����Z�:�3\dߟrN%�9���H�5
yo{k7O�(=8֤�Eo�-s:9�΍��K�!T����@>��ye�V�c��׏���5-�S+[�(Ԟ�%��L��0@x�� ܏mx����-N�Fζ���(���Nr7x��{�t �nY�yɲ�z�N#��ع:I>A�H%]���Ѻ�Uſe�}#c3�K��A���#��O?EO��Ɂ�
�b?��]�ՉM��$�qNzhp�@RP#7�wjwyr2h,MV`��*�3�"S�C2Zd��nJl��	2�S�+���IE���i���ϗ�,K80��a4
������r�F��c��APь2!��#�g!sɶ �)�qnE�`!:���c��aΧ/I�;�˕�4
*��a����x@���z��/�b��x���_�](����������	��U8���b��O��"�ʗk1+R����C�_�m͝�a0�( �]S���EA@N�T��M�]d�0��6�d��T�D��S�}+�6�L�囅�CIt�������J���ذ���z��r�*���*)j��ܢ��ԇ}׈�s/uTd�=���P(g�u,cm���'W�Y�iW���<���NB��
6`��j�!�����UXH��U�Tj��L���&~V�M���9ER�7��7W���Z�V��j�~f\����qGg�G��5��x�������w���r���m����Chp���2�kK��c˝�׆�al�b&<����Lϔ7&� m��n���P,J���k�{�����t�d�ts�ȧu������-/�܂��}^�x%�t�pve�"?%���	�.:m@��R���krbH�I�Ĺ�*SϾl���5+�d����8�4#L ����W���#���$j�9�q�t�~��q\�0����S����r�U�7˦���r��4��$���thtܧ�XO@ 8�, UM� d����_3�=r+=��C���S}�����6"�-�Ip5���I��8cV�`rH�{�"�yU��Y2�l�g!�DS�����*�lEc�-Ci��\xF\�=%��7|<�3����0R�T]����ѹ{��>m<�,)�3���;+$����U\$&z�:��͜p-�'��0�m�*�;�!���j|�Ɋ�8t
�7ѡ"G�V:������>�?R'��I��]Ex�w{M�	:J��2#���X��v��l�~�x'�xc�_��>�kV��Qn�" 9�{|�q�gX;�M�'�D,�m�_sɖ/5�MS��y�~&V��0�����DErΈ���BaE,S[?'��r��tU��C=����}��f�Y��V+��G����9}�HR+F�곸�H�ܪ�̒.5��}v���=�'���Z��i��"Tus���y��[֖�;��5�?j9�Z��ll�{�vH�fi��%�_�mE,��7�Su:nk���
_����a���!�wͰ�.����J�_B3Ce���4�*#���i�� JI�p��'�LC�)���.͡�g=,��/����j1X�4��9��_�G�@��U��aa�P;qp��?4�1��L�g��\��-yC���ڴ;#&Kn�5y�D����qm�X��y�5b���i�Eۿ��1S*��metMB�F��o7�HGf=Q%�>J����ˀ:�dWLW��7`�J��kl>n�(���)&xo�2[���oڿ�τ���8�Pu�uN|���[���3!nf�{��4[[��l�u��{�ֹ�D�Y.�����Nw!���3��L?����E9�qV&j�=��G���_��4`>H������d>Q�4y	XVݤp�ّ/��j��	�q�]��9��ۄA�9��_W�`�>�з�����}n�l&��ӓ�D	�S�1����0K�K�W>:��l��D�p�0��j0v�5�M�D��`�r���U�K�a�l%��h*�Ǎg�+,yF�����,|>��0v�ag�Щ�� �g��.Pn�~�D$V�j�F5>�'��U��M;�2�����`����|baP^���5��q?�l�
!ޛ'���F��Hҏ;�j�m�~�'�r7�ye���B	�(߆Vq��ɪ�
�ߋ���Y����M�Ci�p	�_��EPǰ�I�(3/L�=�a��RS&�s��u�Ѭd�ϓ:��HSJ\���˽/�]]M����B`f�0�6�&�B��[+y���e`��_%��Gao	q���6�	¬�w��p�O2$���ێ#�ZH��>�j�k�C�z�{0�	��XK��uwv�(��� Naʒ":>�5x<6z�hڭ��Ǳ:���=�����yA5�R��G�<�@��Z�\�<���1���MW�&l	��J�6ý؂F��e�)���T�pk��U�=�U��a��2nr@yE6������&��ǀ�߬���$7n߁?��m�A��/�Zݑ�_��D|(���D��52����d�'��&w�7ȢB��5���3���Vr�\��!�B�Q��};��ߒD��T�|­$��=���PȋM�{�s������[���~���UO4ّv��5��O��`��U�)E9�R�wX/rs˺�8����R��v��iwL���7�Ek�~Fh��7�v �@�
�fj���i�hU������ $���Tع��l�,�8wڡ����B��`�b�n/��	����̎<�gˍ/˵LD���"M��"�h|�VYm�t8�T��v	�P�N���x����3����i[;��)���ׄMr��3`O�r�,�Oj�0}�j~Fjw��,P�/Cez�(O��Լ�oP��[@��R������YC���5D�u���|`
������p)�G�54��tBl�_j8���w�Z�)���=J��e���Ic�MH~]�h
�:���1d)~.��Z��V���%��^`��I��/�	��{.�l�nV��
Y��[�ˌ�?�<;��t�.m�dM3�l���^l��v�㋹-��H�F�ա���`&fn�-?�Z�d��+��_5�x��OK���tҞm֑J�~��*ȱD�H5�����~e=���w�V	A���.��BP�1�pH!Z�ŚG�Ey��+GA��^���)A�v|�ѯ�S4ZbG%�J-j�v�qA��A,�"Ӵ����y����;�֓�ZXr�Y�C�a�I�.�t��mʝ�O)v�o 3��pO煋G��nD���MW$��W` ��a:y��X��;��6����`ͱuy��?���NZf��$x�U���J�?hg�`�W�y��l��`]�_'-�Z�E�}�/!7a��&(\�d�6��c�dG�7�M �¿�ο�^�O]�*��ܽ��\	B�1��u���:4���͙�{��S���:'�W+�bE볮g%/����!I=�a�O.���%J�=�ǖq9%(=�̿AB���=�7���c�d]1��{T�U�.��B��G��s2�� L$T��������Tұ7���F,����+!�f���Ƨ�����~]�3��ȫ�pv0�1��J�[(`��-�W#nOU ��^8�N��܈�j�ƿ�+���!._��~(ob7��ߖ�v�Y	}PE�P�c�|���e�
~�>)���k���V�c�Ӧ�W�E�W8��(���y���I��_`MH|}���vk�)��������m_*���0V�
�w:#�1 }�H���)�{UfXG�_fՔ�{;o�r�[�����2�'3P:u"cR.+cT���qְ����_V@�m���ݐ��$��
�#D���C��
�H�t uҲg��?"VD� �+iY&��gE�>,��yz&�ߣ�L�� q�\*�e;�����SR3�a|����s Q���v�´���bOn�3����P�"A�U�i|��3�l����Ւ)�kQ�*i��%�wA8!2)�$���`�͢H�NKMm7������>S8�:o�4�ޱK,�}�/�e�� G-��ֵv�d}h��F�U��l���%�*�臖 ���?$<��YG��\W8A��p�:V�N�$�jݱZ9��~�c���w��4�� 2���H2�6����N1�~�-�]-^�0��A0$�>�(����{#�js���Q��D���b?��^����u�C���c����S� ؓ�)��I���Jqϟ��B�!Yz~�����)`�.v�{{� �F���;vūQݒP@���v+��qZ�ZKef/����A7�'6uB��{�5�h:�@Y�,��H��Z�.w�t���e6x���^�ih2���N�Z;#�2�)�ߜ�)���9������f������Ôt ""	jf��'N�ZK�
��3�t
9I�T���N���@�hhpM&do���[����x��$�ȝ���S�
�����s��Q��<nBh��a��j/���g^ܔh�����	�/uͲ���\ɼ��/���ꩿ�g'��i�t+1��<	KՌ�Z��tE3�Ls�i�P��=e�{:B�z��{Mt=��f�m_R�A}KB������<�5�Գ�F�������܎;T��$@��էJ�K�uX��]\^���g��C�oA,�
#l�ڞh�l=�iW֚(]��I-�K�3X;��|&&ߣpY-��77�w�g���#��{dW`��z��ux�q'PC�*�]�iC�q*�;v��Ӟ3�_^2!���ٔi�v��}�6�8����?P=��M!j_�%�/8�����)��})��+�$��o�	{ϰgS�8)%.<c[i[C.i�c�et�S=}~�jG�ܠ6�.���L��|�kC���<���ǲf;AT�қt��:���f\�~���� �m��E�s�=�d���
��D��꣯H\�m�4�ȸ�?�L�=M?{q�D������L%pu��e�(m�y=�:U
�%��Y�g�[tY�eIF����0�e�ظ�xZ���܋
%���c���> ��1��R晓���7�X���j���;�>���V��k>�������Hw>�f�1*���z�|�+	rp_��I�lUh��?�^��i�Jr]]�:�b�R�܄�b��ܠ��½p�/M(7�Y�:��HD��SLA����x��a()�YT��0/�}�i F:V�4�k�]�A/��#����F�5O8���hА(�����"��pR�4P��p��iwSd߀ ��Ԑ���+u�}���nj�'A{�^_���p�	�a���)2��o��ه��y  4�[,\3�ю3���R��@n7@�?	�~���c�Fy2! �F����T~PRύB�˱�x�eĨp�~"̹���j��f�����H*
�V4v���K�=\!GK�Żg�K�s����cG���U�u���fq)���G���#=u����H�X�X�u�_�Ѐ!��*Wz�::9K�Ċp��lvU��v��(XvC�pRq��Wg$\|)��8�V�!q}Y	pɵ%/K��i�a�#c:��҅1����U�ź��Z�P����P�S0^ş��U:I�Y�B�.wJK	A�X�W�zp/DA��oRU�(r"Z�%��wJ��q�/Q
�1���9�B��-j�i�Rx>Ӎ��,���e��4���a{�JPp�ǣ'�����G��&��=,O�͍>�'�60?wr�h�NE��D�GNP�L �%�P2��{ ���أ_���S|g�&�Yu����v'm$�|���rzQ�	'�x����#HFK���)�5݄�����A��ʨ*���%h����%���n�)���4;	����OM�F�
�S�J��}��?���YQC*����+D4-���	!w�_ub�h\���W9��Jy���\�mI`��>[��+hGmtZ�� 9Zm�c�~#S�	`J���s��xu$
J�C�"-D���vP�2Ԧ��O8.�,�^^f_(�p��KNJd���cU*��哖}gSa�}@�9%*��E�8���m���z,vVo����aO�we�Dh:Qi}���;������L�U��u�c�ZdxT��~O���p���7�̰ϔ!���Xe�s�G�m�t�:b}ϵ�D*��3BlD�0	P!��cB=G� E-��(CRV(K�s9;���l$���9��,A�����m��f���}N�*/؄��e�� ���>��A�L�����i9H9Nb��Os鶤j��'��D0>���tf�Ϊ���[mf������`|}��v!(���t��vb&�^a_���L�I�C]���HO���I� /�?�H�j�e�S��Mm��H��ET��$��BnFg����%�V�;��������V�*���g�[�h��}g��� ��^sF��2Y�*{s쐐��nv�d�JHM�NV�p��B?����`;���25��=e�FJ��ꟼPbY�	y��5SCE�1g���v�2��}F65� IyK(��yh# a����p��F�̈́o�x�o>M}�V �JV��4�Y�,���`�L�#GO�Ių�F��{�1+�R.N���Bd�4��ʟ�계�Pd�)�YT=W	%?E"K��;%�ʡ+&��?T�ZN�|��+[Lj�Q6�EI���#Y��z�6�4K�\���� �!�{5?���F1�\�G�F)���_����-��O�+��f�4q�_�`-K���MB���� $�>�x⒕�:\i�0�Z1�mL�B��Õ��=��碖q��ٴڢ ����m\0�+*�&i#��gx{o���T��n%����og��_ZZ��.�40ba�k#����H��n �Ľ��&�c�D��#�F<�d��o_��(�k�j���e���f �l����Q��ƣ��#��(���[俼t�b0J�PZ�wy��
���iΠ��z���w�X�G!�Y��?�,a�\��Eyh1웑�tkJ�oy�݈fBs;��!�0�AH~�	2t8�+�k[�N��'M�M���Dq�=��:�*��t�gu�B��9V/�ŴS�ƎN��G�PDN%�!~��<�#��_J�@���7����E�AI	я����D�j �ɓ/���2�
�c�=s�ȃ����Vq���e��x;�I͂��b�/��r�Z*(��R�ɾ"��Y�v�>T� �x�SzO��{��Ur���h�7�>�������M(�Y�C��:r�3�MzA�x��7a���u�P�*Ǳ�3����
؍\�����J}RV�����
H�u���p�AsG��G{��xqeW��t�o��d�/�E깜����o+*���4�O����z4\M�uP �G�֟2k ?�ͤ�]$�md{���T�ЛHtf�����a�teV#���*|XW�NfA���Q���MRx�Ƅ7�Ew�U�&�ʨHc��:�ū7�@F�*V����A�U���o�xA�;5�G�l'����R)s�S�ԺC�����q06G�h��2,���;~=a:l�^�Y���{â�Q��Xj����Y��4	7��m���*9�=�%��^&��T� �5�_�L9=�yT��<�b/Lq~�wo)iqO'(p׾m+�#�Gm�i���Ff��O�s�P���ց쟢��8FX?��v��!�qX9[>�&�O:V}��wƧf�Pa���hH��U&T�4��cǿ����A�:�������LR���xJtn��g�+mS�F���XwȻ?T�,(����y��\�SVku�It�=B{�?y���
�}��X�Y��◹0�)b%e�i�7��}���Z���-Al�L_�S$�$�$=�9 sا4���z���>8m2�jX ��|�l��!LMB9�hS� B
�p_4)$���k]�2W[�b��I��Y�v��r,�B=�@��6��jx��Ɇ��/ՠ�ၖbR��Ws#)���ZMŁ����x���q�}"&��x�NA�s�O?#��0��O�ϕ�Q,[�Wpk��#�0�[JN,>�6��S� �F1]׵]�k���%d�w�>.�%��4h�g�4G�6o�lYu�@��c�w�@V�s�I���]��?k���R��UP �iD������{�S�^!,��8�J��{d~۫ l]�x��@ܕY�l#����<L$A�z�����D�'~��׾�X�a*w��vZ�ި���wWUy�'���K��rڽ��:���Q�p�*�B���K�\κ�=��q�9�@��_3f E�Ru�Wm�Bŵ2�Cu�N��h�(���,��VU���X�zJ��1�ݗ,%A忢�K7�0�!\�DB��S�T�1̟�n�(M�Î8�8�1j�' �[tQ���T���n�7�����#���C������U���W���5wYq��Ǩ��x��ζ���Ά�����q`~	
�?�����){��?�X��������@U��^����/K�6:�jj:!���"�a������(�0������&U�"5s!�ޮ[ĕ'�U�FvN���K�N�sfF5�u�G�38�'�j�v��ӌ��5�h|S�Y�]��:-Jf�gS�ۉ�-�;��[�̺�ʤn^�o$��@��*�rw����a<o��h}�8�K�@e��d&�P3W�w��I�w�E�h�lR��XtӋ� �<o�d�0�'�r��6w����PڪhE���:�;��\�)�u��+_�y����Q�{$g�Q��W~���0�-Ka�e���g0ʶ������d�M墀�y��rlF�0M�:�]�1ڡj}S����5��R�_*</21dZV
��+<�l�B��ʍ)W�bV�c��B�=)�c
P���O �S&e��9ՙ�]�^y��҃|6���á��n'}P̑y��L�Ǯ��Ogfw��[�,�o�fY����0 �{ٮ,Yd�O6A��1����.�.��(�Y=�[܍M���i�_��/�s��^%K�����d$�;��O^LqB��EcP[9��z����dv��6T��A�ِ}�;KSvz^���[�8�a�{"6��~�������f��F��\��65Q�G�5|�����+��F5��?jy�Bjo_*e�:����)�
)��i�#����pbOb�"�؆��.��Z�W �v[@��z����M<ܮϸ��� ��k�\�ļR�z�)���^�(V���շx~e���6�9���L�.��S���d��%�S,����b�����ئ�۽#={wG%��Y$a��"��a�V�kҢЕz^=`������b;U��~�Qz K��a|�7����!;�sV�Ň��|�����f�)��
1<�b�>tԜ~�C�k�=�l
��ҟ������\$[вUM�7t�j ��m|p,�s����L��}��u�	�o�e,�y�|�In�C�
5kp�����v�bF�c�$]*��j�"����4��(	M�S�h����JV�Vbms�mˡp���يUuY��'�ަ`��jl%`:L�v褜�1��$�v�+[*e &�z���.�i���i#�_�h㗮"�I�#�CF2��ձ�|��5UC�ǽ;PyEDz�x������ׯ؎�^΅/^�Q'�!���.������p��M	c�<�� ��?�6զ�F��a{���9�yB��.ݖ�nܽ����|�w�Y���wɞ��.r|�������C,��4ծ��ʞ
���<D X ^^��H�*���񭨛C�D�
>����+����=y�c5.h��ҧ�u�X%�L0�@`{�:Rc���U����L�
�	N���s�c$�M�� :�΃۲LS�>�S��9��f.��3&���b��U9s��YL$@	�Qȴ����m��=Ԅ\2,�BB��9g6�?�HV����v�1�#��2�b����$���_�K�"�� _5Ա��1I�P�oA�����̛��ܳ��(2��{�m���mL &�U������-b�l?���w����yH�"��I��j�5Ă%��>I�>̫�KF"���L���(ؐ:�#�֗_I͗V�+A���	�ʺ�+R�F�'��$�n^AH~�.%J�k�t���56��a�<GG��$N�h$%f_x���:0|���6�|����:�?p���j.��
nNp����l5��|�Vh�������傰��/�����6	��N�B�2����m��o�
 À GB�~b��~ٯ+��<�P�P�b֋i˰�U�PT ����Z�BpY��+$s�p�������Uݨ�zt.oqu�4����58���k'��{&�&��ft��%U9M��%�Nf������9YΒظ���r�X�$�j�C[+cӂm��oY%�+���My�[�f��y����Tj�32��q���,'���(VW\Ay+D�؏�\��J�� 2�۵��(QlAѓ%w�p�����3��:�+����ˡ�J]�@@9����@U~W��M4|H�1�:-�@T��"�Ç��x�b7;@lב�U�����H^`��D�f��5P��0m74�q��M��i5����EZ���?}@�=K�=�}A��<s/Td����m�*Q$�Y�.�"���)J|���	��?�-Ĝi2Q��[�-TiU���!��%ӤJ��MT%��oŨi��c��w�q���y��u3u���߷G�;����>|���@&:�j�tKp%)�����N��˞�������;����WD�	�#4	g�z�ڜZ� �����((�8�!�Q��T?��3 �Cqt;p���|~�^͗�j�`��Y�7��{�;#?�r��u\оRċj�*�c@�B�H��_��Tal��`ZZI��X�6|/����N' ��}�i�aN��a�Z�Q�� �����:�9�Fën���|��׷|�w}vƔ9��\�1"@ZH��f����Z��->I�S���[&ͤ�t�\��0`��=^;�~|޲�_:��9��P�j���*sD�A~������Z�;�&Az؆��|f�G��Ρ)i��H���<�7�N������SU�C�U����d~��^Z�@�p���G�v��F��M�L1�<I��[�p |�F��]��j�+�,��4f����ӣ�UA޶)T��%���&�*�8��m=[��!�l�}k�!��d'��f~.��4�p�y��;[�K��L�=�V�6�M:| �`����j�
oS��q-���~x���l,�KK��5�J�Xn��XSܰ��7����,�� N�ke����`%�N=eh�9*�HojBb�'j���x��::"W?n�j��)�ȏ���W�eB/�|$>��$ـ���)��&�*�j�PUk��m,v��Rۑ�̔~&�����ܕ��F$�l�� ��lɔbŝ>6�V���"��L��pj�1e@��W(���v�CԶ�=zڻ�6�hnG-���L\�]uU�����Ay�6�쪿��t~��9��l�sl������:����ZWL3�1��5ogr�qv׬m�x�K9���֐��W�D�A���h�h�RS�ЬVk���6�E����M�'d����Of�Gw���*S�Cx�p^�3���g�O�L���߹~o��%�F3 ���T*���y�؃��� />����k迼�΃Cջ>]�2���x�m'����P�i�oZJ�*��@,o�x�~͐�.t�$Q~'�`hI��>x�?AR����y���.s{f�-^���^�x1l�:,�21�^c��1��	5�%�~s����[����ߣX6Xd�6
��J�����i8X�d�;�!$�6�gZ"�z
{�	B�6e���B��8�~��o����>��|�������u&Tߟ"+l�C�j`�oT�y�a���
^�2�/b��mK_����j�Qj6M1Q���M��F��5��c��@U�Q��=��|޶6I�q�vSHE��B�[�HiVs�݊�6�o���~M��L|��j<,�w�	=GQ���	H��O��Pr���r�$�\�'d:��q.SI��9x_�T||ܐt�"�{-iw�붤�r�ف�%k��^�B��q��B&�)V�y2����N�_�e	�/� -?ŘJ�����h#5���x��d���o�y d���:�y�3/}�i����R�k���xT����l�c�y,�J�o����frĹ��~��g�Q���p+��.����`v],6��H�99&Zv��O�OՉ|�2v<���p!>3&��E��q|x&��Ԋ�%+�%U'�l.:��Ǚg��3mA`_�bz�4� D�ݸd�i���o�W���A�z��<�����U����[{�]?<�̬�1�.}��S��BU׾j��Iσ���!}���������b�7���do�c?ed���� nby��(/R| �UYa/�<�׽"���Y[�F$��� oC�@:r�Ѩ�El��a0�Ŧ���6ޝ�9D��Gr�d*�`x��<}�;&�I�\Z��-�����)t"(%;�r�ڙ��Ӻ�T|t\%�\�pѫ�V#9qD��g��u��s�O9�Y>W7��+Wi�}����Nj���DLآ8�$�s/�N�1z�	2�:5�^�SO�����<I7�'�I�df�M��|_�{jg���~`�?�m<���U��Y3Tf�Ab�'uwλ�;���r��X�,�䗬��ɘ���%�Y:�=��vr:T�`-1�ͮ�!�1-�Kml7����(1�������ڿ��l	��j�MI�"m3����*B�~KS��bFS�6�*D�L=�^�8g��<�7�&�q'�rHx��}�B7�`h��wo���UÂ���M�fV����&�J)=��Z�����+(zUl�̻[O�j�nӳ�!S���{^���ͤ�=���:.��c�|o�6���F}S�T2�d뒫0	�ڿ��s8�ad����O���!@O��!��G�+SI�4řs�7�B�-{����pq�̙	&��t�]#O���tco�Pf����9AϣN�خ������F���@��YY��
G>�E��8 ����k�����B���H��y���A ���e�i�����y8�˝�Q�_���
�J�X]�R���8S3�d	���,ԓ������9�a6�vѲ|��y�O�5}5(dͮ��*�4����jgcJfO֒$iDL� �f�(���iF�����?�:�n�ٸ'�}��V�U7ngɍw� ��p?�I�e)Z�(G�0�N�<X�@�J���6���	)�)P�wEKފђ��%�Bw��ќ/�]R�L�R�y�Q��;��W�2�����A�KN��r��dP{(�bS(E�:��V.f����[���l��/�?O[��m*�t��b���D^��O��`���
����A0�J-cZ�8�<�C� L���rM!����T�� Y�̱{��>
����c�C-7��P�RN'�F�	���ƶ
�*�r�H�XdR'	&ic��R�l������)�M�s_��>��~wE���q�Ü�-��t���(�����n<�x��]��Vh�	1C��ו�j�6r��� �g��+�������nٔ�"�R܀���XE<y2݉�U�A1z�[�;���Tv�d��k�f��� ��!�%KL��B�5@O`q�'D-�1�@t1b�^Cs6b��G\��Fz�㑃 :Y�?�5`��Ȫ�Q�E��۴��E`��q;��֞�R�L6��TuWGK_���Q���3I;�������p���cZNg�|���w�,�W�l�����ZQQ��bտ���BY�"���Xx(�|�R�J�U4Ѕ�� ��
sD�����" Y�ù�ӧ
�W�(zD�?�Yfk�*���*�؃d�_�OlKn�œt�P�?�%�y$⧒�P&w��.�H��ǖW�QxAic��/��>];�(�d��f;B�%�P��=h_& nu��YXl��x�@�3co��V;���@�5��]�e׶@:0��-%��5�eV�`/^C��mS�ȅ�(��w�bm��
k�<M.�̴��? v��>a�ؑ�Շ�L�o҈��徒#BF����������$�?-�>ά�]��ɗ迍�Ff-��>��O�-��Y B�wp�AQ�_���J^�N�Y&�nI���4�u�$�}?8��"���kQ�Q2�'��$/6���:L�D���
��Z��������n�����L-�n�Ԙ�k�nrH	؂ԠJ�I)ՏX<�q�E6:��q���|&���>A"��{WA�U�t�l�k����\[qA�y:)�0a*�[`BU���>�X�$�>]�F��ǰȑ�{"��(��������\�{����y�_�����חͽpҭT��g&F��P������H�tw�D��Zp~uZxb7��4A�>�3���>�)���Q���Gt�5�Գ5�eB�x��B��!��ٯ�=���F<d��M15�������d�:OYΠZ%��uMx@K�Է��ə��Ĉ�x}��⑾�R^�'�ُ�j~����<����k�ص���Dm�z�����T�+.�#����(���Q���&���$Ee�y=��:�F������В�$�@�""m�;LH�>��)
�e�B|M�"���cep.�Q�>�o U
��C����� c��U�)�7Mv�a�jԦ��8���`����+/u���s�ܱ6�%���]_����)`)^AhT��-t�Bj���-[������`!��⻥-��F����\�ڨ�q�/y>�I��«� ���K�X㖳�54��1mK�R^[�u����8�k�N!]�����G˗-�w-�+
9C�/�~�����V�]�����U�q�Gb�����F��H�|�z:��̾G���SG�vq��_0�B�s e�r/��m�Y;XNYoo�z�J���J��y�_Ă�-��!�ʭ_��u38�X�a;�+?�V����	�Щxi�ebTGS�H9�'-c�r��������1��Gҏ(0΄���1�v����)���Y�7�=���@Dn5 C+b��'q�u= ��#�&i[Q��9+�f�׃�n���[��g�V�X�xp{r���D��N�w�&�9~�Ã��d :aS�<�9��]�fkЅ&Y��h��ȏ��fW+�6]iNt9�*��<h���^������%�>�*�()Q}��nq���n)�1��JsF���~�TG#�#ߦ��n��VAq�,nR *_��aeTɘ7OaF}˒u�e�<ԍ]�:��t�.C��/+Z��%�wWE�Q����N(-�+w'��O�\z�U�W���Z��}D���'d��nU��%��7�z6�dl�}<X$��Q&��4j�K���ͺ����]w�u0�oq眠�����(!@��#� ��Ub(��|�w����ղ��i#��{V{_Aq�����r����!��w|�q��)�6�#E�20����К�:��OD�A�d�K�����Z4���T�,w�% 6�����3V~�PoP��h��#M��1FO��}��-��Ѵ�
�W�14-�D��'\d�B)�Ǐ&��"�B�VM�c�����!No�E<od�{���aM�Ae�4m7.�Բ�j�lV��&4�R1��L��?�	���e#��5�Y�k��G�F�I���Ȁ�2���jP�Qn��w�3.ض�d��G	~���-�R
��T4O���Ȓ,���,V�˝y?�۾���zL���%}_��Ո���M��ˢhb��*��\L:�m *&0IX��j��hD�`�^IoKt����\���J�����m0� �~'�h��𑒓$ș�����Z�O��8~���QG����N�]�>���8.Zx	�3~%�Z+�.E���d�#��p��t�Y��S<4���F�>WYR�,���Qj����&N��+Z+�o�Οp�Vэ�޺���A�΂�({����6���ݞ�u�Z�!�T�z"�l�[n�=Wm1X�S���Q�!d�@w+9�LTX����
`��-]e�ȓjyu��j��*���h�*$���3�s�
�*��o�p487���7�� A����,#wbPU#e��=��zB4ٕ�Q�\�k��\�(��J@8X�wOl~W����q�O��F��2��bC��]L�%���V�	�'�Z�4����<�5b����B��2���'�� ��9���T���ň��(S�i�4!=P�G�
.�L�~G�����:�PqI0n ���qݤ�Ϭ��"�蟭l -����W���{0���Y܇����R����+G�W ��K����=gE% ���M^\aB㔩�(}���Y8>��C$>L��R�qS����j��J�R����.�#@Th^e|��kCJ�O�GT\I����9�ˍg���0��!*�?E[��;�ޚE�o#:�=S��PN���A���[�{b�Tc��E*z�F;�ڮT�JG���Q���S��?�`N���3�[@��`h����m��P9-����Z�ZΈ��� �̅�<���� � XT%��M2lwX`Y%KUP���d�]wü�j;.����0�D�U����g4t_���B��� ��j����j �,E��S�d{��H�{���V��^�'Ni����h+�k�8-:���N�k�ze.�e}�#�6-	]����S7�l[d�2j������o�҈n9.A;�{[f H�,]���YR�-�X�]�e��ï������?�Bӗi��W���+B�j�"fM<h�1(�mnGm��+��ֳ�������Lp�Ȓt,��w��兕@��Z<��'�cp����;�v}���BXd����-�l�l�V񃧡�RY�����A�[Q*��P7/���"��;$8Bؼ#��s!��Ck��S#��8���_@��
U���4�w�<P�w��S/�Q�2����{��A:�����ͣ�g��ߌ&d,�~=�3s��jv����f�Q�؇�c�%���\V5����;QP��!�tb����?xyj7��*Y�4�X_�r̠��^�� 4��`����\Xe[{eO$��'�܁�s�9����Ȫ�].�;e��8]5�����ϵ
'-3�1�E�������	�i�b>��d�^�͈���sqL��lSs���_0�Q�B�٢@���_҈�p��,�ad
��Ȩ�X��"D0w��W��] �0�y�p,D"��6���bc������ߚ><��ȴ���M;'d��m�%I? �pAM���ܐ}?7�c*Y�*������n\�[�t{�a�E��*�4�*�`�}���w��T�E�r�(>�(��1�0�p����ϧ�5}u�ewmcK�+?�����PY&�m>��P�)�5B��Ȓ��u��3.%�m��Ȑ��B�F����{���>:}Un�-x�V��Fh�`�bb���E�Uڿ�b=?�2ym;H�4៚?��l�sY��Y�J6U�Hy�sQ�� ��wC�~)R�y�L`r�y��q�]�Xlb|�*��-��~���Q/bg��S�}5��Cv�{�5��>����3�=���4'��Kf+�J)d�hf.Q�xe���
���v�s;�'*1DJ��(���=�;�P�j|^�>!L3�ɶ�v��z����"�18A�1��� ���b���WY�}��\ ��ߎ|r"#��N���1����%n@F�CMOm��s�V%Ŀ�^(���㗚D6u+��I��GEZ�b����1`���V�I)��t��a�Z2��̗��ө-�Gj?���)�|�a�j���g匈F?��#t��-�ZF��iB�����gW<�e��v�� �>T�:F=���m5qb	�V�>�ŧ�h��MT���}��#��\yNR�)-�10��t�)� "O�4
I��G�L��
��tD��q$k�?��-O���/syh���9F�v�$�2��/�S���[ԫ�iq9����l]��Ւ�� d��zьE?�u��wy��9���&��Z����IG=ˌ�����xK�'K�҄6�m��b�	3�r��E�{���S	�����wLo�fJ9�&v��㼞h��9�w�mAu֍(,��}�V<^�`�ʴ���<I���>�1~H�~خ�y0�Y��_!WYO���J����k�̅l��F�'���}㞝Z�$��ɕ�7E�Ke?'_��bqG�.�����ln{+-���s���S�U�����%pD��(��9���_#�X��QWx�� x�"E�νL3[��)H���C�=�Y���r�C�S��]����R��
X�Ëv���
�U�OPm�lpo�yE����go��3I`�4z��+B �U`dEQ�亜-�V�[�.h�P�F��`��8R��R�	��S���w�OK�=��-���h,���H�p��%�6�͸嚯&���:b�/��s]n�ۮ������/���XO �$�*e)�/n�
�~��
 ��7�����Q�׸��2�N��8Ƃ��Ak6�I;KfnyI{�S9O�%�}.$�]����.�ƞ2�*V��R'�OT�Lcq��P�fy��Y8Q〲��*�����mZ6�8f��e�GM.~p��?]â&�"�G��nv-]=+���c��nn������$$�+dw��r�!�J* �	^�Ī���]yH��F+�]��N�@@�h�iÿ.�v�.�\��V�T�k��<�f^���Ng�N1�<,5�0����o�X�+�:wi�~���Ur-�vy��R�L�:URL��/��	|k·Q�F����^Ě(��z�W�����2�3X� �[�e�D��]�X�R�#��\��d��]_Ȧ�;N�10�Xs�L<��4I�v@� ��Qevx���c�t�e,2eX�#��� �����GZ߲[�hZFY�vTJUk��_��U>ei�|p��!�d��EkN��L)���{2$�sg\�u��-&mE�	�[(a�֢
�vj����2�
'n��8Lf�JE�A��V폤ᚠ`2/������X`�ht�a8��y�A>F�P�v�˽��������I�3.{N���z��a��#�X����=�N~�_�J7�M����k}��=��}u�x�2�͆����D=��^�l�sEu�!;���?6�΀8<�l���d≧ �7�P}�Φ]�{P3s�[p���F�D6�_���h8B�4���I^�C9�7k��"��)rt�6
��r��}巹�T�M�]Xd�H4���d{�(N�'V)L��S1cn��h�/!�1�,L�ѕ��tCA_�>�?�(	أ�ϝ}ZK�Z0ݫWE��e���UG�q���!��G�΅����>�I�3S�o¿O��zb%Y��w�tlzv��n!�E�/����v٘l�	T���w��r���Gv'����xN e�bv��Y���ii�����z���u�ܜU��aqqaI�T>w՚�- ��|�I2>S˦z��,[n�������o��M~��M�5|��x=+]���'lYs,( H�O9ym�[�W>������& @.tj��A	�?�퇎I��yz��ιŮ'w?��a���PT(�޻�#D"�}#Y��7�qg��X�XzӁ�C�v��5,�@/���6i�����\�NS����=Թ!��{�����
��[mֱ�,�����u8��\u�6Ig�n�@��q���9N�h���\���c��7��&�G�ĝn��������P�c���ʴ��j����B�&E�шe�R.j	��[�iV��u�Cw�x;��C�'mbM�of�=�UidB��ʺV�i�7���9ۄ�kkW�$��$�~��c֊�Hp��<:n*5HZ~Q�w8l�C���X ��U��LϏ�]�B�HQ�o����T����E��Q�����4W�D�]�׎�IYcn��"�K@��ߴ�a$lK��Z��:`Mm��_ �H��FH��tչ+�]X��__�6����Vۂg2�����-����^�/D���׫,{+G�җ��R�ti�(pI;i�X��E�paOn��Ћ,�z�,������S����w�dT�S�<0��2�^�,��1m ݓ8�./��0j����x�|A4��ܬ�� �g�~�৻5V� � ���bF���~�^C^7/�}v����h�������4>�`tV���Oh4�r,��f������Q���ߐ`����t������ ��hLTI�+��{**� �S��\�GŔ�!s��a�A��Ը�I��Kߧ�t_l���l��f?:r�t-s�4�}wi���ej窋�������,-���8%��n�"*��zF�� ��-f)lj��>a��d���ްj�N�)�K��Ǆr�b�����m"��z u�
�Q��H���)ة�����'U�{ة˻�О���=OkT�ZR�re䰜p꼌p��)(�á}�N��<�Z">���F�sk�nE����Ⰼ�"�"��	�'	z[ʏ��ŉ�*�6w���U"*�ڜa�6мx	`�۷ ,����B��;��1^I�XW!����7 ɚ�A<����BM���?y�^��>0nW��ڇ:ɢe��D��J��e)$���ѵ��p�3��#Iv\ٛLX��薆���g_D�.K�J�~Ч0.s����ϗ�':�ɞ<�XeDz�=�|�ap�5G����.	;�d��ڮ!�D�Z�u�N�J:~��m�nS� c߄̱>+�=*�R{-�:+x\�6)�t ���з���x�'�)�A(�c}����c^@�~�`<�b���?8�޽��s����"�zPF�&�ѩI��XjO���uk�x	n�"�-U�:���`_����"R���f��9�9TYqǧҗ-Z��)N�X����,��SfjR�S>�M��ê�Z�2-D<x�����Ɩ��'qM��i���l:#^XD�aNKL<oz4����O����H���a¬��C�!�����<a~��d5�>6���b�1%p}���+�|δ�2����e��.t��1�M/D�-���Ipd�<�)H��F�0/�����KU�`]N�X�s����0�����ǈ;,w��ݮ���,��i��8�SZ��^�س������cP�����\�es��Cgp�$3F��u����A�N�.|�i��ۑ���0 ! JaYb���:�p}T)�Q�������/)���}DĒ� 5dJ{����0�c�xW�����z��k/}l��L����
�s~"��sZ4�"���T������<�#E��FM�s���|G�"ma�[�w���dA[�m6������j(�����z}-<AZ�P
?1����5@{���T�`����4;n�Ji����צ>G�E.=�h�:�K������V��j*kWħ�V����:L���qǔ������:������h�b���,	c����h� �	��<���ú_�$�{���5i���҆,����m+R  �����}^^�Q�5C��O��X�w��-S�6��?�@����	�\
����=���u�*N�~�Stt��d���X��*	ş��s�R�Jf�Q�G�-���0'�&���W%b��J�z�{�_BCѿ6@���G�����y�����˩�q�8���d�m<ȩ�ZDm$=Ἑŵ�!�(�F���h$/fV�al"��5(n���/�_��:wѳ�"3Yaf��L<�ti��w�Uj�@=PvK%�a<��#r�B�{R��S �?��8�	M(�9_%�}��ˤC�7c�'���Sn�q�F
�P������e+�G��Y�~r�e�]I���ӈ(Հ��6�"\���yu�G*��� ���}��� {7٠��[X����#�6�ԏ[U�6yH�����k����Z�m�=�y���j-DN�F��.��?��i�P�1g�4$j�P����-���;�J¤KEܛ��e�)��_Ԋ""N�u�$9��M�X���a�Cs���x���X��~њ%�y�}�@�ɧ�.��,q/�',���"�dj����1]�i�qFʲF>o�f�Q��ʅ�n�|���#T}/��f�16u!����Ԟ�I+i�0^1��S6˰��C�U5�o�����ښC![ץǒ��Np�0؋�9?u,�Zhj��J }�A!��D�����0��C�����mQ.���Fn.D�QԮ�QZ-`���rҼ7?�[�H��}��!f� !�"���];9�h� z��7�~�\p_|#0��7}1�*�,ކ�����8���$
;���2y�)l��&��7ؾa��/x�`��U`YR�M�{�cE�[s;��W�q��`@�wu�Lkぞ��lT��K����¥�V=\PEZ�S���c�S^5*U����H��6N�;�%A����a��*;�?�!�v�M6J�k� �E�%&)��W:���g�)�E�B�ʟ/�-f��1���iA��k�z����HЩ��B�����$���W�y���g��*��Bc^ϕd�G�c�+�ޕq$������j�2*�N�o��l�WR�;�ft�[Y��h�B�#�zr��t�W*� ���^��#*LZ�@��cO���n�Ɏ�������̂��A�KÇ��!��lf�C͖C����V��>�W"�����	�ޜ��ȹvz(O�hS8R��[�o��y��آ4%�ow�cV���_$��h���'7�����/U(�����e�L 2�)�V�A�!e�,��e��
�0&��=��9hdܡ�&�J=��L�.;��>���{"`)����O�giKj��T(����T��VzK"o��q�U:�
;9�ټK\�dz,@V��7��r��wQǌ�u'wy ��+~�.^�����
������g�cDW�d�ȕ����iCX2FD�9��5'r�U��YO��Vf��О����Jd+q�E��p�N(&/�O�^!h��{����J�7� �b��F{��ٽ��Qw�e
Wk����p�����;�e}����3��B��G��`G�6�Ky���©!|�����&�)5�V�k���i>�vC+�(�� ��En(�ŕ���<��e���%��Yg�-R�m�nԖ���������7��:p�O���x���G����:��/OkG�+-:
��œ��?အ<Z.�ך͹�E��!��;�\�ڿ&�m�S���;���b ���i�^щj���W\MM,�B}����ƈ9�eV����R��ܔ�?I�������l����FU�f�^<�rQҀl�S�I���/jR5�����j���P�������������2vb���=]��Ð���d���5B��v����/����C�Fǉ=��G���?�GZπ��{_���"����C�d��=)�2h\�b�d u9s�£��!sGG�\=����8�P@3�ƧË��\�NՇ��<���}���KY7�5�Cs�"�^k�LuP�٫^w���X����k���0��-o�6��O�sm5GZ�4��Ƀ"(a���Ү�O��߾���i��w�2�i�l
��bѻ��Ao��:��,b�- Sc�"�WG~�u:��x�wg۳>�K>X}R��&��؏�]*qC��@�Qʛy�*ԇߪ�>���yH���$3������"E�x��aX�h�@�\���� 0'�X�p-'>����SM��	=�b�T�+b��'з�P>��go��Mݯ'E8�B�5%�S� <vDz���l{>_��=~d�1̋)hW��y���!�C��i�����j�,RU����o�Ћ��ć����QA��S�l{���h��X��2�?&LK������ՙӭ��� 21�0�&7g�Z$+:P	=�$}h-E0=���� ��A#?�fF#��6�ҝ�R�8����U�t�5�VR}�%zt�X*H'/컯���/�w$���=�_��
 � �'���c�t7��x�@ˮm�S�g��$
8��V�&�g	�������r*E�W��Gn��|+�%��W�	B��+���	ԛ��{^!�n���ԚTg���~ �M�����D�2��Y�pR��ȍ�{E�� ��>=[_��d��14s35�`�C�`���W�>�.���e�	k,�L��Q���D9%�-0w�5l�魎�:�S����dML���E�/q]V
��4yG�jY:�\��DGT������n3�^E��zD�|�?u񏙗kQ�����WZL���ʱ��c�ف�3��~�����zfkR틢�rzz!z��#�%]����j�lʞ�O4IS	v�?�@�k����D�L�r�KP&�_h�W�@������9bp��B��y~yX��&������Y��D�V����*հG��#��)����A�-��J����'ɚU)�]�H��=�!������������N���\qL�)����X�N4��w��>����I쓸#7�a�����"3�-h���N� &4�R��؄I4M��u{��z�l�Նx=1���҉q�Th�| ~QH@�?RY���n�\*�Py)ջ�e�8����62%U �, �iC:E�[��C�)����L�\<�g����]ޒ�`���ԁSB;��K��z+�A��ѭܰ�,>X/����f�bԷ$m!@һ����:�z���E��w�H��y*�J��Sα]��R�?C�=C�>?�X�d��#�	u�Dᆥ�%��o��;�v���	`����8.�L��4�2�)c�!�?�D�;�[�eB ߉�#xԯҁ�*��׉��gʎsoQ�ֱ���}�-X׌u������`��>�}џb6�m����Pd�0�� ��L�n��8:+v��)�o�����`Y���o�8C�;�4܏R�6�G���8���sf�>ц����-H��r�d���k�� k�9�H�D,�v����>O���]c��x|"����\�@)h+T�IcT�T�)ӹ���y]��Ҹ)ܐ�ܟs�������k�d���J���t
=�<��*1UvK3�C�*���t���X�a��{n�S{�^���L��L�گ���;~��k�b,��R:�,I�h�u������E���:��GGz�A�M�łB�~o{�1�w�0pEg��[?��E�ʥ�yj`mB�Eɛ���Ұ���͙�DUf�8{X���'�Q<����"(�hO��g�#pg��T���d�6;�G���͖1�I��'�GťG��~���	<���v�6�i_��Ҡ��×*�yc��g���l�\:�$��u�T�޶� =��S�D�<��av��Ī�7$-HZѯ�:�:�,�c>�6�=hs�}%ߴ��nJK����Aho�+V]���O�J�N�%ꯁ�g�`B�V0h�x��������@(���5�k)Ce4����<�6Q ��G�'�>ӵ��#�1D�z�p�>�׆pm�?E��'��Ǐ��J�9&Ÿl���5+������ۣw��9�����q@��M�fo�:�e۹�F�AU��k���;�$ �fׯx,s�%����i��h*M�䡍�׈��K�5x��Y��	g/i�-��V����ֶ��jV�^�Х��Ƈ�ʽ�m�7��=ZT����wA��ѭ��+L�I~-�n�ċ>�܄�*��[��0b|E���Z���3�������M�O�)�%�m��Ժ�ܵm3�}�T�P�j<?"�H/3��΁p��������W����ۼ�3��\�f�C�RȂ�<(�Z�^Q3�oo����(�鷠�2V6�n�<t��t0�`�cO��ѧ�Y@������C���sw��\���\?dZe��i��͠�)�6|XG�vMl%`�5R$W���9m%J�)���r�`��dƑ�+ۅg�{z"�ǎ�3=�3�
�E7�I��f�nN[߅-���A�F7�O��z2�yiNxxjx��A���Ė���V��&��m1��؟6�>oW��jK<���,v����3���4���h�p`���<�쪑~�y�`0F�I�j��F*li%VR���-�%�B7A�r��z�'1�ܜpX�V�E�W1�ed>�!?��0��Q�ц՘��MTYnQ-��\C�^�g\��J��A��\��W'��~�h宆�<�$�h�n��Ӥ�n[PJ2��K�q�s2)��_�A2˭�c�����}{�/�آ*�1d#1�pt*Nkա*B�T
��������h�*#7��%z7�zر ��G��1��3����tZ�y9e^�R:-�4����@`��@�F�����Ӭ�G�)�54Y#��=([�G�l�㿕�}J4.r���X�f�bVH��9X��{�4��%O�f�c���_��P��R��F#xᡚ}�:S��֛Q@ :v��>w�j�bX����GF�Ń�C^���z�
r�ao�I:�X��������ʾ�d�J�W�QG�Y����~e�h�O@LG�ޗ��&����}��J�rZ����"n�ձ�g�R����n�5�E̿�i�Z=���<����?3���cs:���?]���V^�����4(r���Y�x�}F��L��\���v�˶�c�����e�}�e��f�����5�	��jDʉ��#uZ/"8c�>��  ܊�BnX�f\�����춮%��\F\�E��+n��������y,��c>O�%��;�'�����q��M��u�������M�Q���{�]��ž�B�����-N����£,h�Cj��_�wl'�M&<�g*'v{��!��3� ��@M�X��5����m^��92:Q�n���F����k��{ڨ�x���9јd�KB�7�
Zsk;;E+�~q�"�ڵ�0��� ����fq&�Ъ+D��M	�ȣ*���l���������k��7X�(
b~"���׷_3���\�U�)b-���*`+y����l
rHp$R���+�8<�{��Q�&f�_�rc2�e���|�^.M3
ʭ�C��<���o-��*�)`�6/L�8�+����X'����������>���\
�I��,��?ͤ��B'�8�˗�Ӆ,���3/V����o����ބ�d>�yMKaN\��D~g;t����/�ڦ�zA~��O��	���$u���2���u\6��
н!O.�u茂;�ΦX�͙�G#��Tl��s��.���~*������O��Ɩ �l�����ٖH�p+U@��g��d�����D(�E��p�oE+'GL"��C��Ttm�N���R�L���#0L��LKׁ�{����������
��:�Ήy��:!�Vs��,��{�`��V��n^�}�fL�Q�xa������7KM�Q.������:�p�f'�G>��Կ��_�k�X�Q�[wr�F�/�)��|47U��k��\�:�9�fմ�GN�P�{�+'�f�v��y)�ȭ�3�F�ϩ+M|�4���)0�,�<����Z*�޻�4h;u\�t�V'�:��{�����H��������N;#��#����B4Ȥ���Z����ܺ��������H.�SSt���=%��{WB�V������8 ����հd��D$�u�������L��V�kO�M�0^t��t�^�qjRZ�ͥ��!$��*�����$���Xl�b7!S�\بb���F��yל%�5=io��Rs�G��r����0��������1��2/h�N��wbw����L8;�/��2�	�P��z��5o]otVݧ�|��'ܨ�M��6sk,?� �O:'���026[͓^���U�RO�պ��K8c�»��"�.��|��Ѹ��/���!�;�EQ�B~..9�i����0D�������.Bru��/;���d�aL��~���]^!��7D�(%�w��{
%v�-Xs�Ƭj�Ǿ,w�%e�#^�s��dw�d�1�ydڕ�>C����)p ����K����!(�E�Q༺I����������L���
o��o���m氝���Gj�u����́�I�^8�.�?Z�����ŧ�v���qd��j�d�y���G$-2�5��[���Q��A�Ү���(�	��j�?��阖2����������8�c
?��V�W �$'�j>Y�юXy�£I�Іo���UX � �O�;5��<��-P� ~����
(F��T�R�C�B�k��(�A�
ͽC���u7W��x�Cw e��'=!?9�&�����|]��7_�0�͖�u2��ٶ��I�j �p�#�έ32t�x7����#S6|��6��1�	��]�;��:������|����	���P@���P�hՋ��?Xh"�'W^�vу�ؗ��X'��<���U?UYSp�=��v0��|����
� �	o3�Hw�K
�<�T�����'!+y9I��$(�ӏ�.����D� �9���+QC�}gD|q�}�zS
�M���+n�����K�Mz� �?�������(�=�0�ӒT�S,������� a�]�;���2G�_��4�d��b@�� i7�J���Ac�W>R�&=v�2[gC�	�z�~�ű���+�(�C�%�H�o� ��'vڈ{\I�7��e$W�	]��	�1o;��-��s3�4�.+�j�o�����@o���P�ܷ���'a-���,8��`�⾆^U)���=7��ϵq�W����2����TT��!~A��;~� 1�@.�:7ك7V��v�2�:N8��;+4�f�s!=��-z�[�\[+ ��������3��� %r�j[����]�6�|�Z�Dq�e��c8�/��8L���cEMӄ���C���Ǔ��/�l�`�ػ/��(88AX��}�22�����1� ���a��В@*���>�Q<���s�͇����\O�-V�_��3�	(�c 7[�5P��X$Z[���&h���ȥJτ��� � ^���0i��������/Pπ�#�s��0��&��h���&��x2qQ�_È��mB��`��
XtR��0�ˏ��������d~d��"�iR�$I��W�R-�ot���_�9?F���:M;r��a@G�Oz���f�b?���+�4�io�>�m����9V���pɛ��������I�g���pm�˅�L=7<Sߜ�]��%QW�P�Eo,��I��ߔ�U���V�y�(�`YQ��y��s��s�h�FK�3�S�Tk�[\d>����f��Ux�Q�����3��_��l�wyϩ]�/�A���k�wt�������`�p{%�{#3�
{�f&�����.ӮU��څ�\��58��E������]G6$E:C8H.�\+Kp�N�9Y�.f��Tk*�R���#� �sۂZ������U}���m���-��S����_g���d4���[P�"o��ƿ�x\;��8�%�	N�̱P��膷%H���o��� >�[�u�D$LK;]Rv��%�0�Gob�]�`dv�G3�lوp_��E���Бb��B�|{�t��)0{`��U���RN{�O[�l�ɀݝ>%׋�z!(0��0�ɩ?��~����\:l�=OW'�fN�	�@��.�/7>��T��H�K�z�u1R��ug���0�����!O��VRӴ��.��TRa�*�B�޽�Ѽ�'�f��.x��AC���2�o �=�4DJ����H�+t|����}�	6�^^':�M�>_;���Er��vJ������H�!f��}m���M��ū�S��f�zK$�_���>2����&c\���>�L�i�76�jr���Jl�]�F��a��%Eq����#��������2�����̥Q(����e��߳��gB]�F���|��(��Lh�I$s/�=(����+(�TY_4������Jn@u���f^+8�b���ާ��Gg!�e�^�w��>���įhLrmY,�0��G�($.�d��s�;�0���6'�uS���n��y��y{�f1��`���I3�+���rO�yE����(�qgC<La)@a�����X�L����;���|grʌ$j�,���s��\�	Ԕ�H<�-����>�]��b��s�]���ocS�KE�;��t!p����h�R�ػM���F�0�_��f�� Lp-$*|�y`p��L�(��>�Ⱥb@%��d����a+��:�Y��x34������������� �<��]�ܞDT�kp��u@(R?��}�|���m���.��l�Y�Į���P�Q=���-��Y��a�Ο��O�^�����kth9aV�$��}Vo�g�X���_�]_�l"c����+�F5n+=�������%��h���'`��-��tKx�$�,��?������aa<��u"�祩0/�9��e�J��٠:k��J��F��\��
 ��pX�s6@�����[_1x�w��v��?�h.�H�4��A �ߞo}ԋ
d(�I��:�r���$�o���e�ɂ��|�
4l�����M �a[�O܀qHd�� �_�R���Ƒ��%�A��ݯ����~�Pbs�$��ռM�D�]t� 7�U��^�O�M><;?xcBo�e�s�>�w�ܓ�sk$��c) �1�KXo@`/�YIH�V�3GR�����Z��λ�E?�=�����x=�6�	�*P�y��8����Pf2��T�!�9A�1��T�uTM���n0s�63xͅ	gB�Jp�NB�@d\��$�S�˖�$�kW)5�����ݚ��KyYB�?f�g�V�s��]m�e&���J@ή@��-�>}lDJ|=	m����t�۫s��ĸn��� s���0�P�b��VDޔ=^�+�Ed��,RdP,�'�)�n�q�"�4b5��G`Jyь��RE��\r���7�*G��1z�a{Dļ꾧�_�ֲ�X�m����Ȏ��zG��[� ���������!4�	|����8�h��i`v{?���x�jEŨ��u�4#̔�����CZ�`̠O6'L�6o��@F5�h�իk�9�´]�0����0�fU��q2F�4��Af���#��v(UP��e�f�6dV�����}�>B��wTr�h��������!���qBW�Ɵ�q�RЇ�"�n���|Tٝ,�2�Jm4�}�NId�ș�Np�j�LN"��a{��(�t!�E�$���p�.�#+2N�D�o�Ύ9'9�a+ѡ �N��*��緭v�3ȵ��菣`����h���^G(�| 2(���.���Ə�Tg�)�h�y��, $	��+��O䯱��*������x��G�k|Y&��N���}�g��^����N�ڕ.�)v�
(��8����o	0���a��l���0��?�U����L����a�2�@�j p\_Ɩd�ޯ�ڟRz߿�������~���ӝ���U��Dr�cw�VX���������#��b�sY֥�� a;f�f����m�p���������?	���D��׸
?��G˨@�K�$���v+mgƋ�Hj��'9��9�ZRl�|�"JM%22�5��y�ɹ��f�Uy��U��7�編�$Q�?א��:�3�0"��b��P�Jy:�+u��֪ߞ"�'d������g�jN?�c���ۨ�hTZe](��BT����F�{A?N���;�~l3��h��(��BŊ懮^Nf�'l���2��Y�吅�lA���,N��k������ruh%�-s��^4rg�
�!��8�Ή��QH�\�=3���/����zqD�:֫�Pǒ[O	z��2���{�dw|�5��s�:�FLqM��qJXUe=lh�lC�DH��<�e�Ժ�q����:d6J��Lzq��eC�C�_�S
P;�<�����)�ʳcl�JFM�On��y&wgTlhH�E��hgi�`oz�K�7���H�PQ8;�:@��ɗ+6����CZj�в�㮦M���U+.6�o����X���X�(Q�nٌ�e^�eTٷ�E�-�����k�@BJ���3t������%����O~�t�"pn�1EMU��W��r;�S	gԣ ;���Df���m��i��8i��� [#��탓Q9wА�v��]�{D��㒡�U#i����ua1!����[�-���F�r�i�C2V/���?���h��C�Kc��B�!}1�{�(rB��}0�Їܖ��͋�p/���+*0t,�$@�����\̶��,Ѩ�h��,��	m8��zuR���c�T���u��'B)(�j>��������kZ}��C�9�M�5�5p���O{<������$�v���	��*.����Xx��C4BPa�G�,�i^������h�sqʪ�35�w;�e�;K�Puj*׾5.� 1|Ag$�Ҹw��'P��%T���>[�S�}�T� T�{�����td[�;�s���c~�Lݠ#��0�ɝs?��L��įbH`<�AÙtD�+�����c��Bv��7�DR����=]�5X�k�Z���7H��/���k���i
�Ix�^���*�i�r� ��A���fNK���=�`gߵ�\�@f
etIͶ�I7faI��q�4qh/�|(�J��D��]�f��ew!�ڎ���CE�u�Aa	Aƶ���U�3��APA~;�d��Cҁ��8<��cN[���=�]k��k��J��x����>����$K��u��?k���)	ظ��X��?���YsA�%M#�$=缧���(��ZP����+/���Y>�pέ�?0ݪ��\�_h_�}K2q�ߐFX�U���� <웚��Q��O<�##���A�$��=;�J��'Ҽ���K-�л�z��:���ca���ٞ�G�P���}�N��2�ѻ���� �g�� ���4�oR4��������%��=3�.UZ��E�h�I�!��Q��>���{]0���6
��tr6��U3q	���N2�ш���n�}���@����4q;H��*��n�7g� Pi4�]�g�7ܝ0ߗ�~v-�Bô_���oMc�C�o)2�0}ӫ��ǿ{��:��&��}V�_u��%}q>��t�}���iP���#]�d��N8_�Tx�	=�$�T���E��eIY�?����Ow���f��g��2�y?�f��ꛂ7��א6�2*
�#%䟮9�{��!��E���춵w���(�V��l1-j��̃��%eB�9� �/����Y	��UJo��� |G����� @�\�%�9�y�G�s��_���ڿ]򏧔�}�0��I�%�(��`0$�ރg�i�Fx�6�E���}��T%�1�:��l?��i/Q���*W�/U?�|�D�kN �A�1x�-�� C�b t��]{�%7݅��]cLro}��Q�R��}hR�[ɲK����lS"y��J�p�乐�͂�#��N��Z���@4�=�����X�U�U��%U��ˮ�1��@���P�qN��+��CX���7 �4 4�;��5Y:�6���ה�B�{=�p�ϊ�̀�x����8+7ѴZ�a�����[�"�,Jz�%We���d�zk$^Մ�|���Ϸ�B_!1��m_��0ĺd0��t�¦w'�rl35���1�
;����1��vO,q�Un׼���:P�d����;Y�Gov���.w�/1ӌ�Z�%��{�"֕W����#�2�[��|U2bo'dM�$��z=lmXÛ���;d�L�X�o���CL��~��U.�]u,�T�3z[4�l	���T��-(zFLCN�&�f$����y�Br��Mh�faqk�y\���5L��6r�	A�]��OOP����P���	h������>0�j�ci��/������{E	������Гս�xA����r2��[ ��U�GS)��.���g�ٚx�ū�ܔ��E�(|�{� \��ہ�p���f�%� �i�|��[�f5$o�W�͡vlZ�6��D3��P������A�y�Q��'�V�e��]x��\���!�CwKO!Z�T9�{�矵`-L���>ƫRٷqů�A_i;��GKt�\z5�y��gQ�%\-�o�d�Ԡ�"��f5=G����|#$RW��[�Z�M�a��DFV�͜�N�]=�L�C��,x�l����3_��[�y��s�I[�b��z�F�}D���MQ��!s�pG^�9_��i�ר8j�%l_���	m�Ο"�o��h�z}o��0�uJ[�x�<g�ؼ`k-h'���%r1І�g���~N!ǖrսUKIu=�Ӭ����<����:M���@�[����{	���D�A��Aëd �ͩ��`{t7 jz|\�T��]�'�r�+������<�c�:�Y^ O�������[��3V���`�ҭ&�5�<�!7�:S>lݠ��){r�'�Y긖��}�x�R~b-�S"�s��8�h��I2!�F
�GdZ"��*�0 ���P�S���Y��IpsW���J�܊�.����
9 �<����A��|g�ZI�̍��;�*��8�p;+����/�LEЮ�P|=RH�vU!��:.#l^+�+��d�'~7xy��nh(�A��*������o�H�%�?�b�_gf�d�?���ɨ��)�]�\]���S��˫�p���R��� ��D�`�V��r!ק1��pZ�g��9iP����ʄ;i��``P�'^��%�6:R��8�k����ǭ����9�À�ja7�VE�$��_d��s2�cK�� �X � ���[��?��a�����Ӟ��4 ���R���o������a+� W+�_����O�k6=���� �-�	����IꏁZ?�᭟$�Amm�j����u������'FId��V�@�De^�j'-�i���daq�F9�o�_�DU ��}�-���|Ȇ(�h�k�
�rx�˚SY~0j�zsĴ6�[�$�}Q����|gi'�E`6�<�>D�EW"�b؋���j]u1{bj�T���lD|��C.�\Њ[JOJ�1�w���;��,����AE��H`��
1�����q��R
������ߔ���2�k��_%)Mq�b-���x��åBk�_�k/�.P9vt4{M2�V���7!2��-����
:��pPgyW[�j��-�|�p�������,��R�VgWx����:���} ��H��^ӉnZ��pI!@ɝ|3���\.������86�m[��ύ��QH�������}Ӯ;3j�R
���:�����4�@�I./�nƩw�97����ĝr%O�6���f��;~ېڃ<���'��g�ne��g>��.ai�G�n��]��v�؟��ad�&ޠ�9��P.;���,�D k�#���]Ą X�(1�R�/���)�`��X�^]w�$b���k�}k�	�L�ͻd0�G���u��D�X���~�4��|������ަ'�$��C9�A��
O�5%�bo�٨ǯt������3�:V�7��i�}�U��2�U�S��X�W�v����<�f�H��� =��X~�ǔFK�C'�ř�N[�(��Ӻ1C�4�!CF|;Β5lBk_�Gj�n��������Ë�E�Ȍ`jBC�F�^���	�~: �o��q'G�������f~��\�8Y�������E]�,Uʩ��/$�n^i��[v���R������$!kt+�����,�SL�Wv��E���c�ۇp��`�*~�V�c���|4�1�p}��0����	���L~��e�r�)ٚ��L�<v�{0>~/314l�x�@)qA�$�V_�jUȕr�#-*�����fL���q >�:S�]��H�0��@�����t�	!��.��ϗ���iI������×Q�=�K����7E��5� ����%Ⴣ�f~9`�R�G�>��p�	��m���N�����X�JJM�NBaMiی��㡢� ̘J�d�G�����ݙ�Ն�{�BʂT��G�i}#j��۝!%C)�v@�-�\���d�鵶v��G�e�C`���xY�IQx���]"m�L�u�ǎƲ�7M�$�{%x����T�	`"��(!a�3[�������'�β �桻4;�u���;��ݭ�icz9���3-��l!�e�p����Z��$��������TsjG,2�r��x(O(g� I�u,.���N:vD���[e���I'rf!Ȉ�C��-%"fg[���Y e;U����_�if�	Z���9�����#����؞A�q'���]�*�u�F���#��t��W���?xT��l0U@�Ϥω�1]�)�J\mf��f�O��0��w�=D�q�qr|��~qw�����1�S�����@�D^�a�h�޷qJAXYum��l��O��FK�_fl�����k�=�AV�ْҠ��v��!����<���K{�S�<�	B�v��f�覵u����I@�u�4��QYK؂ ��'���й��^�܇�1@G�:t�cf�aua�%��Ip��u�ץ�>��Ur2O�(5���	������H�N҈G�^K��G��6N!=\#��?�%
��ʙ*K�beee"�	��-�?,�cK�v�=���q�RN��f�� #<�'�x��z�v�f:l�k�u�b���
"79�n���gOO���K䓵9V�!�M�2�U�`�6j5��V-���K���xgM�ۮ2l�~����UV���J�5 �'ZM�bn��=/1SR_h�=d�+K�3u��#��(�U<XԴ�d����p��ٚ�ܖ����!÷�
�r��t�����Y�v����0<�{�}w���_���\3�U��|�����e�`T,���C�nyGT��n+���~?3m���K,�5��U����>�G�|V=4/h�8����a�h�q]_�ȟz݁
-�A�;�\1a���=r��N��b��Oߗ�ov�Z��Ӟi�\4���\��d���>�S������!��S#�xOk�K��CeJj�"9����c��g���!f�cE*Ĉ�2����&�^D���M%��h. N1哆#������؋�ow�����+�,_UJV2_|/ I�''!^4pP�N�!L��g]��^c�8�zyל��Vd�ʩ�?���X�#��B�����I�_2��d6�7F�����&���1i?�2P�M&_�S#^�`I�d�#��Q�^�Ў"�N�w\�Ŭn���z;�����J��9�R��~���}�ݏ�������r�+�(Gv��^R�1����a�J[0��UV�"%
d�k��y��}�Oa"�j6OC�[���O�{$�41	�c^�V��'bx���٠HO�9X+�OA��}�s³��S�F�X��cȨ~Lg5��E��D'9zIx�C����Q�-0:ݪ�$�Ш�a��̘�s���� �d�d̡�슦�1��-����!V.) E�B���`�@LhZ�ň�� ��܂7]��r��ǘ6�U�~��ނIf^*aQe1w�č�y�yZ�-L�p�i�Ӛ�49,�YdH�,<<GklT����X��O�r|+>�V/��"ܛ�m+�hv���ͨf�j�q��>�o"�Al=\�%����D�!��=��7O��CL|�o�x?�n����U		� U*&2
k{��B�ix��)�F+��l�@9^�z5�|��
]x�m�ѣ����5)̃��i�~&�IVuc�귞?
�}� |(��եzn��d����/�ц�����!�@�n�t9�<tk��٨�� 4�B��9�Zȃ�t!�I�k����3�����HF���`�<�v�םk9�]nfv��/ك1'�=�� �]�	_�Λq��[�g� ق�`���2RO��_,����?ܾS��hgY�/砷һ[˱�Mt�W�9�������p�v�o'ZRJ��O�>!�p}�i�&Pv�qP�X):��w�ܳ9|����7����Լ�ד��14+�޻ִ΢��"�Ԡ]?�.ȁ<� ����6����o*Ob̈���7rzͥ2��ӴY�Kyx@��E�Gv�%R=��p���zϦ��[8���l0D��L=O���PdZ��KK���c9\d�Kyquc��~8dsT4�$ʼ�Y��>��A�'d�
��wi(�K��`���;�/���Ȓ�+1V'�ﷰ�;9���MzZch�E҂�"vըR�q/���0q��l��WR񿽱b�Y��Y��K�H�jE�R��U�	sF\���u�I�ݶ�#-g�W2F�'�靑�?�G,��x,V�T��g�Σ���V��θ�-�Hm.w��@K��!����w���B�X�RS��d�c� 3��;d�,ЪPɼlݱr�ޑ�Zw��K.�I��P���Q�������@�q�>=p��(��f��ț�o�{�;R���̭IM��qe��/rQJ�`��$#p��Uf:`��bk���3���r*#^`a�I�(�O�J�z׃����r�E�D�g�И�9����֌�����h���!�u�l��?R�ġEc�?t� �K��l�v`�6��UP]S[�U}#���������b1�č��Or\�r���A#��o���	+��|��E���*��"������$�>�+x� �j�_�>޻t�����>�1�'���,�m4���pX4�@f�j�%{;�SLa��Lܾ_�󄑳�+�D^�;G@'R�!�a����m�{���f����������Ep������X���I�Ӆ���}Y��!�j�d�Z�Ǿb�4���"V[�k[��8��5TNao�
�+6ǔ�A;��=i̿�ܝmƓ^�H���y��s�g��f�'���(��-]��&.�
���W�N�A�}o+�R����_�be�s8�'�:�C>�P�mZ�F(�ڇ�RG�[Km��JJS{��y�����B@�w����)y�����8�Yʬ|y�ǀ�V��Lg�5�Y�L���`���3@�*}��^�JרQ;��ڜ�/2e�xjc�5�U���of��;��Y�p��/��v�ƀ��� Z�,�د9�q�V*k�\��Z�ٿ�[}��Ц�Bg���DR�� ΁V���?��k`�{9�d��W?��+���a�E�c�����M����'m6�����6����+L!į��ǣ���	/q��UG�ϻ6X�s�A��B�#¹m�	�����s!Y�������:$�,�����4"	��֤X?)��.l�ݹd�ru�@O����,�}���@���)-�� +L�(8��?A��ee��w�����ݛOW�T���H��,���y\�z�w^s����K��f%�Y�2l�A�H��ޤ��8
��8��%�ހL���#����K��SY�J�����-y����vY�L�WCt��06F0���t*�-�� ���w+�3f�Ɨ���Y�H_i�� AZH,Q{ɹ�t;�tņL�=���g�~���r5Ў�s�]��n��e�8�wV�F�{RZO�ިQD7h ��3�Qϑ���碽�0��A �h��$	��0�C]8�K�l�h2�5K���DT"@dp�ӫ{6�??7u(���F��ҰR�x�����PM�ـ�x�3���R=�Yp�/)�/ ��r0h�@-܈�1g���T��mZ�H�B�������Ef�p�!%��bY�e��SQ��y)��2���r�WL1�u�F���"��Hig���Sھ��(Q}@F�����6�6����#�s�M��(`������~
�`X�[�F���*�ПNm�!V�e�7Һ�)����AlȽ�W�:<��R-�HC��>�72O�����I�융 &��Ӿ'��#v�3�Mx�N�7�V|��j ��D״\F�N�~P{ 
N��,�<],��F3ߛ.��m��p���������v@�}����*1��n��h����]:�a��V�j�4ng���Ck�O�IU���ǚH-�ïAi��9��`-�n|���ј��2����P��s�z.��)WY?�sU����6�n�Eick��P���?*փK���}=��l��Mbr�L|VY��ɛ�z�`��h8�����D�>�����3m�q�Qj5���M�90�3�
f�R7�	�=>�ta2}�lDY�0����,��6}��?�M�o��ذ���u�Q>��Pdn�S��j6צ�����Y�fvB�B�'��(P2�f���[Hu�VP�|�KSV���+�E�e�.[0}fs��W�.��B�T�_���� �|�Y.OО�9�����e
)׾Umu�]��~�D1�n}������>�x�nk6�X�@�m�:�`jl=������3V���L����#��B��ŷM�5&I4����0�/m��<�#�}/���+g�s�pJ���i����~�i/�#&qU芓��0��f�2��'c��E.�K2MP�)�����bi?c���N
�x���O�}&��Q�%@ϿXo�*�4��������Uf�HΫ�]*���'Ҥ�!��ei�`�>����ux"A��RWł/죊^S!egI='=ۅjP>9�ܪ�M��r��A�˽��P�J	т�.i����"
�:��jj
\���v��ٔ����h��7uBw�ᝂGR�q����)����\���I���?u�)��7���+�o(5�e$����6��*F��Xk��y���)�֙�e)UW�yz�3z5˒VO|G#E�t�� O*rq�U=i"Ҫ�!�+���9�ׁ)u@;�{��A�
!�_:;nTz�뛚ho�~�[Ȍ��:�d�bK�^0�7��"ʠK�>̋�.W�.Е&;H�U:�c�����I#)>�^/�Z#����5!҅[(i��qu
�H�??�?�=�|��5�2'"�4z���}B/�
����Uw�9.����擂mu����R����A�W3�����4���>���7uq�Ԑo�-}nf�{s�0�t��a���#&3W̞���H����R8s_(�?Zl�ճ���S*L;��%��|>��igl	�;c�������\<��N�Ĕ��C&�jQc+�#���sDff�B����']$,󁄚`1�W>H!+��e�1ɒZ���Ԭ��͝�,����<��e�:�e2��̭Q*y3�	VvV�}"X�q�8z��E�͈VtQ�i��sg(!y\AX�rf���UK%h���օ��R�C^/�عXZ��)�N��/t$��a��4��M�ڸ6!�V��hT����Cgȃ ��#�YO�EӾ�U���ת�QW	V�>jW
�[_@��=O�Di�;�U���et.G�������k��-ʅ��~��m�[dTI��w���}tҾ=��K^7����-wrZ~�>wX0�_T����qL�xj� �s�-�?��7l�z�0o�i����r*�dg�yZEbn����8ld�����Mw���|�6����^�(Y�v2����|��܏��O\hd0��:T��>��j����q�m(�ѻ�� �8\A���*�A����m��pƇyoR���,��>�t���?�l{�6<r�~���wlPaI�u���nq�Y{l|�Յ;�2��䰩�?��[M�4y���:���Xr�#�r��t�hL�ixV��:{��V���2q�c���̔��T��Zk�I�;Ɓ�d$�<sAt Ib]��z�`6-ш��<ΒE�t��S�ˁ�/�[�30�se(�ep� �Y ,Xq��\�`�2{1��}�!�K�(#���3h���G����1����O+��TE-��S[Ԫ|W-�@�lvLedV%5�(9"0�W�:ckӢG�L|�9�:\Ht�'�����`
5�5?�n�G|�~�1~��r�,������%ֳ*��r�,�\K��c�Ե(&�2�:�Hlo�}�	 X�1����ܱ
3'��6��Bf*5G��������Cz��I���>*�?�L�I���cVE�њ�����b&��#��c~))b,;�@�4stl��{��&�ս��7�M�����os�~a^�y��b���U���L�"Է	e����N�����0U��	�C�kt��{�k��C��^aC���baQ߻x��@kg�u>�s���N�ەY4��ֵ�o���C�;��{��Ŋ�����!;W=��K�|6�w)��E|��!3/t�`���<{<N���3Ozr�#��箘P�4uN�oS�������������܏ل}t/��!��s �q���~ܧDjy³����} ���8�>ve�)�e)��D��	7a������;��,
���e�B+�\�����uW�2<���M{�]Ǉ���(�P� P@!9��\?����QT�^�ꃍ�(2�j&�lK��[��duV�q�DWm)�S5�S����4
�Hl��%l��ͼ���� ����d�ۿ�\���%FI+��z``aw�>����T�1X��?��MR��j��kk��yLM�q'a�����1E[-��n>�X��e����Lh�-\�g䗒_���P����o�}�=t��_�g����(��CL�*�$T�T��6�#��������Y���ZzB�&��p� H)3�$�p���_�<[�W,�f�ξ�/�,vi�h�E�Zg��&E���b�_;;�Y��>x�t������o
zgƯ��Hk�Mv�KA�@���t-j���J���ж���f}3�>�<5Q����C�oY����P:���Jzf@�bn���@7� S`�l���1s� �����o|f����Z��EX��#Rr^!{�u$"����
ׄ�	2�%�c��2?�[�+�d�k틟�H��ߛ�W�Y9�l��c@�;R��q]
iE�����8E�en�?@�B�^	����KK�3���yi����+���7���<[���#K�e��m���g��Lٻ�{�I�L?�`��� yW�2��
߂�j�/E�v�7�急�.��4D��XJC�LĳmO�uJ�l��-���@f.�O���9I�F�&f��"�ӊ�90�om��� �S�٤�= �fobX��_
�+wA�Y�����"aV��F�Q+=���z4��ג��P&,Z�����.��<�4�&�Kt�M�����2���>GC�HTd��b׫���X�����/��}��P�O�׈�A(����ܿ��^6��]�Qqk"���Г4]���$[Q?��o�X2��@	���(�~"kvV#����/�!�[r@�*��,xuT��s��y%����������K�E��������<�B�J]���e�`~������={�g+T��0.1 _~ה��M��
ޙ�=6.v��\�ּ�{���_�2b&��-�sn�Qƅ3�F�6MO��M̋�d��3��W��,yͳ	��:�F:k���p��;(��f�JB]'/�=:�Z���/��+8uӺ�!÷ƿK���@���n�5�=$�r�z@��ޓe�R�N٤�'ީ���r�g~I��ŵ���p,M"t��j���1��i���nf��_�r��8+\V��k��3?=�K�$�����d���D�qӎ�����P�_�0��[Y�[UUj� p�}3[<0�MH���{M���B��[�F����$�Z/�Y�=^vۺO
�{����#��{Z������ړ��wd6AY.	� �8�������N�{��XR(>Q[���_�qT�ğbѽ��aGd�BX�6D�诨�x_T�V��\v�@��2��bm64\���SQ�X�oV�̕��#�J!f�!�7������D+.lƀzŗD�x�X�D^�Xrw/l:���!#J��Ɩ�%z:LY:�8z�h� �����P��B�Oc�[^�jw80�*���/}�ª��Fb/��멁��!�``x�������zc9z�Kw�^'qɲ-F���
Q�8��3�����/ptJ V��Qz?z�(x �Pe	wxL]9�~��E�Q��\�ێ�J�Ȝ�E&�u�*IBՓ`��eEJ�|�Ye�D�[��sւ	L����3�K4V8S��.��I�%s�u{"Z�k�O���K�2��g�|Ң�d�TO�E~L��%$Բ��f��"�ŽM���[I��1[ji��" iW�_=jcJ�82)��E�����S�x�i"�����S��ȼg��>hN!���PCE�S�v��Н�F�2ą�P7k�
��͆��=������j��
Q�.5<((�:�9Y�l���`zRh��$����'>�ؐn��9V���z���)�%zf��
�tP��$��P�H��?
��Kb�n���3ȣ��nE��
��Ҫ�S�;ȭ̱��ٶ���:��	�@�!�7e��*g���X6�v��Ybܴ��Ml%��%v�4:��(�j("�{�q����@�=�.�R+C>;4�cM�֡��wDl25��.�qD_*ߝ�F�{�l�4ŕ\U{�*��I�OF5몟��	M�"��m��3d���J]� 5�\���p�W-�����dTt��@V����rH@��(т���W2I��d1���q����R2��W�1��su�$�������B7�i�3!�ÀKz�����>�}р���<�[h������?�X&�����5pQ׻/^���irI��w!78��y��OT&��Če6u0��8r&����Ҳk��}�lP"�ŉ��&�"C�܈m@<2�=���ڌ���>k���R���A��7�Z �{z�2;(�����w�`��	ơiD2�h����GW�?�����!��쀆���Ɓ�<���'�뛒jp 7�[�G�� ���R{�H���G����Ԁ��k?'̗o��ɡ���KU�j\�݋�_�K�$�b[�&<��#x_;�BG��m�����1=�H&�b>;��
W�+��q_1gB�Ex4*�Q��.���J�wȂ���6u<yr����RA�(y��x�e�C`�y�(NO��Jݦ�	�=?B�ż�@O��@Y������R2Δ:�R�Ɋ�}ȃ�VG�^�����sl�����j1r۹OqFv��̨{i��'8]�ӵ(��خ�h|��6J[8�ФFҷi�QZ%n?�v�L�j�͉�ߞ`p�W���uy�7�̂�[�����6#�EN4�ʅ{��[�E>r�=69�k���Tx>q��,L�����z����ف�EVGN*F~���&�	p�%z���U��PV����gf���Pkt�}��(Ұ�L���1ؾ-�c�6M袜E+�@!<	1!Z��X��lx��M���I^3Dv�}�ķ��M�$j��ɺ[ƅ-Z�]��]��aH��}��Xu���w�$w�H%��� h������
[��r�B���ߘI:��_5��t	�D5E���W�u�Ę,��Ю6�<ýi�����h���|Xo��k��E�vS���3.Pq��J&��(�m{=�s��kL�N Y��_���~t7��N�v5E���ʶ�v"e3'�K�s���Ts)*�F����[J�=�%{=����=��E�챪����h����I�C��<�cG�R`${YM�>z4*�a�W�<#��Y	s1�3���.�gE�|;s�4�w�N� �.�җӑ���k�B��2�>m������F��2;���\͜{�g���Z�ڻ�>�.0Z�=zq4����;��.����3��X��bx��&S�Zϓ���p[�t�z��_�
��~��U�~�����rȓ���;\I�1㒑�2�v���E��r[h�hԙ�dn���P�X��|��+���'���A�t�l^in[��ZtM�B�"$he�eq�Z2�r�t��D�)�"q���ܳ��\�@�]@���k#'Lش�#��k{� �J�������d�=�{��R]����B�ϥ�o4x�ܐ�p���[$��R�J�2��~c,/&;���,Q��~?��rԜjuY^��B���$5!w���U��
��HXƏv�3��GY�
�|t��lo�[7X]=�������(���T�ݵ8,�U-��~�,���>����Հ���U�x�a���� �5�05�4W��8�#}��4�oeoЩ�|�%_aM�X*�9P_�>(i��?��o$C��O���14y�O���]/�.�cDl}1rѠ5��N���>�w����U�ț<��h:�HQ�c�|���g.��m��.�����w�v���7mܤ�Xp���4G�,��fߨ'�����d���UL9�G���mt�l�g�6BX�[���T^l�R�>a�s&�v���
u魲h~�O����A�-a�X�(��R4���f�]��C�z�DZfC_L?�k�~{�d�$�+?���0ò9}��,�컩�A�p
������ZzF[m]y�С���E�������bt�T�(��E6,㹜o�8 �2"�_� ��o���9jde@����-UI�_W��3��=�f<�F�JR,6єbԟ��,QC1}��&��ߕ��B0����N��2<<sh[]�YD�G�~�>ϛW Y�9�e};�zB�#�["	$����Z3�>`7۶뤊�i<������f����-���+��VDGV�������W��n�.
�R���Nbǘؙ�Y-'{�n��^吴]V!� �������%���6�+�SQ5����G��%K� Y�jK�ފ7~�k�y�>'�>�"y�Lsn/<N���xz�٦)���/��5qDk��`�������ƾ{���$x1��2�F�ѱZ�u�EV�3�	)b�X>&*<����ts��.ݟe��ِ�R� 
�2v~�c���멯i��
�輒o�	��o_$3��{��Tv�k�^#�`ޢ�,,nՂlHh�t�:3+�ek���}�S���G�վR��ʪ�a�,�F�,A���4�yC��� w�6f{�Qc����� F���$�Q����W5�?xسn���(�-c��1�^���-�A�q~�A?��H�������jYAΆё����>WH�m�O��ds�ZQ���I�����J�`dw�Y,�\U��<'����=Us�6la()��w��A&�z)�����������يT���(�uX�4Υ��?�wO��C�m@��պ���L'^�� \8�c�7��N�����!'�]e�q�^�������t����'�e�"�^J<����ڤ�Gވ�2��wYH��cl�
6����t�%��]Ԝm�A�_F�>}s��Y-� p���L@�~����3��=_�p�1��ش�9q��]PCj��A%���$J'���Ȅ�8pr����+>R�x�ha5�y�-���/��u��N���5rќ�ܴ���x}qЮ���$tk���=�WML�����40bȐ0�z�X	��^�Sʪj���5�f������e�h��a���a�0z-�;�����?���t��:A�V'�Ӡyg��}/
�гG����Sj���q�@��A�	���U���L+�&^��R���=�W���EJ�q]S��~`W#�k�$C��m~hWqP\��!�� M�!P$�6n%f�
�tE�O���I��O�0�s]��j������ŏ6�Siv����X��U��z��W�$��m�§I����2�Y�����׻	e=���<�����2���}T}�L�������7���!ն>��B7���*�i���l����_��F�{�����S��W�WY)@�r�FgUw�]woK��#N:�x����s��Z*����Y;g�P;�F�Wgv50ړ������h�wl��l� �t5셭����W��grv�՝�<y�)(_	Q'����>�!�@eO�w�d���D�<�x���=@XE���:%o�E甼t��8f�5ɯ����B���,�������؃f���@E��d�m�N��(NYx>������ʁ��6y�@f����$_|FB˔��C$g���M#n�u	  ��l#�d�S�M_��"G�?[P-d�����@rɴ(��-��o�Ae�Ӆ�r��Y1��|u"���xX�1�����%J�py₆1�����ñ�����(�r('��4AS��
tָ4q��])��6��:. \K�e-T�m����q)s� V{�b�$ؾ<�����=X���c�;���}�qج��yy��"��9����K3�;TL]I��!�Qp���\\��@��4&�\z~��+�k��}0:)�������x�h�!�
>��UH����;�[�$�[��)j�fjicT��K�fj�3����0͟n������s�Hz�u[8)��_,�[�\�Ț��ـ+&�K��v��꺺6̂�Z����w x1l� a���%'�3,/�A�o΍���lH�u�E�}t
������Vb܆ܽ��<t9G��*��ƙc���M�&��O�5'(���!+��-�p���k������v�y��,�R�H����v����^݅1oAP�7֊�y.�	-認,���G�u��C����8����=��w��(}~4�����h���m��K�rͣ&3�sRV�ũ�6&�`Tlgw>��X�^="�>U��+�Ux���E�FS�u�J�(��fa9"x�����������
�R��Тm�Я'��(�Bc�tX�~���A'������e��o���zx���E�a^�����γY��H���n��ݩ�;+;�b��:��(��d�k�/��(P��5�muoQ<����q����
�t%@�(Ww�V�r��?��Z��	��_l.�_i@J�O�
�|�EN� ���[�/��a)�����%�����`pz%b1~�|J�7f��s^���G�xsf����*t��Љ�)y�i���
�w�Ay9o��j	�}�E��ZVYq������:��w��Lִ�N�����l�st�-^(��VuRͽ��,�3�K�n{"�:�n��@0{=t�5�0�3��|vq���CKԈ��Цl��i�{ $��l1X�yo+0r�_�$-��D�����6�B��2>�UD�z��c���~��ÁW��:A=�N�)��D��A�rO#�L������-�����2�^@�hf,v���h���_6�,�r��8��s����<t�ڹ�I�;A� ��ʁ�������h0�.6�5�g�o�d��m.��sd��RS�#�|���3�$�a��6����m,�CC�}�i~G��L�0z�����?��a�ơ����/ j(p,��]�s0�b,�j�,�e�&�T�NiOevu��r�x��m������gu����Ԗ)��Ux~�nz'2
П��X5�E�<��m�_���h�R�;Ki8� :��Z��p�E���I�����\+W&l�f+�J�1����F��nQ��<ѱE�y�V�7�#q&�q�z�4	ML��{�ʪy�(������aH�Vi}4v?�)T�-\��]�Q�&�� �G�-��i�F��1H	�?�;�=!�G���>�:��`�����Ѥq�O��C�Y@�U$�4�3l��혲�ED���M�ce*[��vm-�#[A:>aj����	j&@Lv�q0��n�m99+��&Aϲ��o�e�x���t �I�}���۞�Ƚ�Y1�]���������.u�9+wY-wW�D t��ߢ���S�����%�l{U�U�g��
JiPIQ�x�A)G*ze0$�&ga���#0�m�4�٥@������������f�� ��OM"7GP�k��e�}h�%��0���sIs��Gnr"�j�ڊ����e_�a�i�$|L�C&z�}�j�GJ!���~v��D��F7�thC u��d�i���ePN�4V�#�s�$�|�'.�����i�X�by�
�����N2����F/!8neb
ja����M��0�J����%��	�6R�:��z������$a� �h�؀A�
:�z�f��_*����G#*>ǋM�j�V�\���Hw�S1����$�y���h������ ���^M�5l�pq=�}���aM��4ן�U"�V�t����\y(x�$������?ƱћQ~ � ���&���)��c8�����(`�h�)���N'�q�)sU�����XG/t�O}Tͱ'U�|SH�F��0#����nd���Ht�k9�%�$f��-5r�&L����o�Z3>G��z#��o���o��6�(��B@�����f��Xs�g\�G����~�+���ч���[2T��Ir��\)o�џ ~�К������ɂ7����R1��rMB!��3H,'�e��{����]M��\h����̫G�堿�ʞ����k��=áͭ�u��� �@���H#�Pz4�о�s�x-y���v�t�b,��W:�"
v�qkB&��m�s?J2k���ƛ�o��U���}�|<H������/5��-�X�wa�h���X̺�,��[8�okqo@��
rOR��R����4us����%|�;�����q=Qw��_y1�(r��N cͳ�!˘��~B��Q���K�k�����w���SU
B����<Td?�>�(�Й���
����k}du7*�4��cr9R,F�Aj��T�"����I�Ԡm�"����7��Xd�3����_�4	��!�,y�!<��L���X=���5Q5���i��U�\�n>'�r��t���QcE-�x�^��)Z�m;�)�}��@CQ����gX���Q�_��`���4�/�lw��I�W�پ��׬�>�SO2�"�/;m��@y�6��MLEI|��BR�\�}O-H��wn0j&���d*w��!"~��1����I
�u�o��yq�$�vP����xRf�7���ѻ�`�f	�)��BzW�w���R�E.�S��=ᛳ{[�:*�����B'j!(�zN!����أ���]d^���rT+��_�袂E������9+�U���_PPJ��}T���J��J��?�׍�f��`�ʲ��Y@��@}����;�WX��~���{Hҩ �"�[Yt�p^u��v/�������]��V�f�^r����͜GW)���<�UE�B8WN��-E-bqU��v5Lg����S(�Qbݿ��q4�uT�;���bxZ�-*����oF�);>����A�J��5*j��p���w��X@3d�N� ?�B�SC��d��0���̭�b����A;��4�<M���c2��FԼ=A�W�Q ؖ�k8X��\u>�K�
q�p��.�-�L�D;����2Lm����.0Q���_�P�s�`� �z�S�Y.�����}�*Uۆ�
3LF!t����-��D�3�'�qcPo&�U�/Q�~���qP��2W�8��ȗ��eNmN�_�O.Dv�
cp��Ev�Mm��g4�;d�U�M�(�db�o����E��$�0��5&��\[���9�==���ť�{�*�L�Ys��ٺ��(N�0�g����gz^��d�Ul��3�4�6 N[�v��0�n�D�	�� [�Xh�q�4��pYu(���f�ShS"<c�ݷc�RJ1�~r9�~�ϗ?`��Bs�!�v�!֛�Ε {�_���!��[&�v'���7�K�jS;���4�X@��$�7,t<)�X��"k��WU�qk5އ:^�T.5/z��{�e�&�`&��W����o������	)�b�ҕ��Fy�f&NX�ɍ�|�B�B\��c���Vi�r���4��m����Ki�['��6�ݓ�I}����y��?���.���f����Ms�Ef�O��ڸЊ-NЩ �t�]��T^��C85��/	�d��Rr��3&�bm�,-��`�X�Sv�á�6"�j
�r7
��d�Q]Wӄ��� o岈e�a��o��1q�gl�r$ ���޼��d�f~�~��������Hn��f��U��qcM���YK?�o�'��-��v?�����"e�?E�q�:�_����=����e䶼<�_h��>(�ǌd8��� �~:�!�\cO"s
X�=RB��"�x�n�c��eG!��+|���+k�-���Q�.9r4
j�'��S���%T�-y�	�(�g��w	�%�k��2�Q7����-��ŴX��y�VB�é�0������A=<�:(I��m�}�[��Y��#b�����(]�F0��Kb�5�?�o|r�J�W�c�����(/�]��L�ɓ Alq� $-�\�}�7�O�|tӪMo0	�X�D�%d.��n����\o���'� �T�]eE�^8��+�r�?#�j�d���`��bj�x���ijPDJ�xe��*�$�vK��W(5\���؊C=����p]]�s�ހ��=W����htT�h�Xu�\d,�_f���J'�;��,�	�\Ö��p[un�n�[����Q�}�qH��e�p�S%��d}������-�����?�=Q@+&MkQ9&�x�[3��b�6�X�*�D 6��!�x7���2d�kp}* !�t�ܳ��kf#��â�E�L"aL�-ò �Oz+�A��}��5�U'܁z���)���O���K��f�TY���6 ��x�o��<X�I�S�O��%{q�6p�Q[W_)����p�ƌ�|IЄ5���e����͝wkB�:fo[uy+�����b��#��0/hmE �R3+���9<��+_�ϴmؙ�3\�MHnQ�\���������g�c�V�i���1�ޜ��&���^��d>�����m5\�U2�f�UJH�z��2�Y�ƜZF�D�Q��z>�)E�Š_~ح���[�^԰o��Pe'����zއ���>Z�>M��7fSK�N-$OW��LGG�r(�<�ħ����BX���g��0�:jH���K��!b��M�11�%����#��5x?��N�C����
�7j�Z�9�A�u� ��GH����~��Y��*`�7������������J���A���h`2��C��;�h�4�zX���C=�M��NU�?��_�w��][#�7-����O�[���β��p��q�ԯ���F�a���q�s;�l(��	�޳@ĥ�r� �=��TVpɆ{b��k����C��k��C��,D�7�"�ψI���ō��£���*��a�f�W͡�����0��Ya<�vZ��=�����%��	d�O`؀�������n�������/��2}�T��֍_�0J�*���5s�r�,�Q�LlO�lg���O��H�ǌ��η����u�Y&f/v+W"ű�*�U���ꭘI�0L�+�Z�ۆB�0 ԃ{ýע��ĩs9�j<�4a&�*�������-�e��.t=o�l� ٺhh�x5kw�jB����w0n�	�J)㈁�!pz�~�+���I����;�����N1z��W�)�i�I�"D3 ��c�R�H�_��l�-����p�]�\s@���xtJ�!0DO`���	|�{����e=ca�*�f�O���=�/�H�xSZ"ws81����q�;�~'��v�BY!f!�dGM�0fGw�)c
�֊~�9/85A��p�
�6�3�Ψ���t$��	(����t$a+NM�?޳p�����tp��4Mm��7�s��i1I2�oN�a�� &�$zd��h�>�a;[I�Ɣ���lź�NJR��1�g����X�1_Mg��rb���Fr���+�3k��ݿ�4�&�owp�s?z@yv8�}�4�wB7���Ձé9��_�J^51�������ˀ�ѵa�Q�Մ.VO�xw��G�?S���"H=4g�5U���Oa�p\���r�c��A�k[k)6��A{<���|�?�79r#��{c�o�ʜF����T7�3_�R��*��՜D��*b]�T��_,K�]D����%+�JK��O���`$-�(b�Dr���d3�����L7����|ö�3�W�����wp��+��ӎ9U���yV�M�l,��Pl��I(m�����q|��N�_�5 L�.��_<%���j��)�b�x�ܴ�2��߯���*!1|+e�@�݄�mx���6��7��E��煽�T�]8�<�9-�S�j��=�u;���F��<�;J/V�j,V��ABOw�0�/���i�R�����@�Aε5m��S07����lq��,\��E]R���o�$�\�d�K���}��t:�J�沣�_ -��&�O�}eN��e�����k&�>����\�I,�^��j�H��)��e*ѱ�E}|;Y�;׶z;&U�~͘��zbB'Yѥh���_���3�	{����f֡h��P�*nE d�2�hn�ڗn$/6G�v�S;��ȐV����j���ÖX��Q�j�Ք��2���=CԤ�y%F���d�.�iZQ��Y:b8�\}��3AX��Xh�v��\a�����T;Ό)\�n��VȂ�Vw=P�3qa�c@
��(�!=u��D��sy±,S���	
���B,Amԓ�<v�GW�q��'��v���7�J��Q�HA8�����U�����c��j`o�6�y�_�1I�㚫�ni���x�,����,�uT��n�&�w¬��6��pFZ�,�m1����D򹕱,�zw������e�!�����kͮ�#�G�i����/KG�g�7�7���h����8�D����ii�Z��9����E�D$��1"Q k�g!j2?�fZ�Y��x�)f����Tz+?�3�7�x����*�����Ӕ\0.�0�!/>���P�_J�e`�RA�򶥦9�]��5���+2��D��ĕ�/Q�m0��G0O�O���>�NC	�f߰ݣ�-���bk�@�2�ָ(u���ms��^%P�����D� ��L8�}W4��I�Ցj�.��\*$���Q~��9�O��8뱰H-EKa�×��
�E�Ē+��m��hn���X�8���`�t�M�5�H�q=�6���I��3�U�M
�Ŋ?M��kk2u6�2Y�������ʷ~y*Ż1�_�0C-J����R����IY�vrE4�yp�ޯ	s؏>�B?���ox頩]������^O�"�Ǐ�mI��9�ʅΛMAul���`�M�ŃJ�OI��j��h7�]I��{[�ew��Q�ʑ���;����R}��k;4���ĵ�s]8�W�rW�98L�2�o��r2�qc>�E�#�A�(�����P�����	������_P0��"4���ʙ��Du�+K��zhR���3ڄ���U(�{#��(�I�/�K���l�P��';½=#����'h�a��qD�cD4v*�8!²�'l�:�2I1p)/k����%k������9@MI���"�w/^�R�]��r]��
���C����K&Hkb
y��JV �6u~y?A(�Hu�q(
���,INg*�Vł�ϟ3HM�hn���+��\����K���S���7x�~���6\��ϵ�\�[Of�i܏�+Ǻ�X��'��]�}�:��W�s$[��4]4�Wd*�Cq����A���b�eH!g��$f��꤉�_��U�'��Q��
��8�[ѯ��I2�ʉ�Z��nHbVzD�'�)1��D����E�c����L����ګ���U��^��� ��]��
�"uJX�Ti�!�W��RZr="#-M��e�Ͳ���E��̯%:!me`�Ղo� Ĺ���N@M�D�ª=��@K܌5���=
��a��*����@�.-WΪ�n�&1����^�X<�r:W.��7Ҝ|_�4C���v�3� ~�RgJTJ<�2�a�l�#e�� <Ȁg�a}w��P!Z�P�<��
�O�a�=5���FD�r���ȑ�����B��?��P�R�{�l�u���yRdw����f ���J������!�k�C�� 0,�B��wQ9�S�<���Z:�\=E�t�s	T�> ���:�&��v��Cs}��:]����}z�%�NP��C��tE��$�i����|<H>��e���`���z7ط��&>j���6v�H�a��H:���ś��Oa2i�)�qa���� ��o��^��ѓtG,�C^Yr��d�Q.ţ�s���V���N�D�\�<.�ޘ�U�uW��R�#�Z���ȹ%�^�آ�,a���z�|.�oF�(A.��$lHE-2*3�2M���Ӟz��X����o��cf!T�%v\Td���m�/�=͵�G��6R�'R@DCk�[�8�<@���X���.�'�XX�w7��(��e��XI��η���_.��@y���g�8i*AO z7o�#����?�p���}~���-5��g�Sp̢����K�,jcb,|�S�Nf����=�D�B\`�9X�X�e��oA���UȖ~����*s#�/Uķ�K���^��JA���<��jFN������J1d4�Ac9rq�?�%N�_Q�s������!o��i��B�s��{UZ�Ϋ06�T�:�)[�'
JV0��У�����6ᣀ���W�5?��}�>�t�>?��JqH!# �{m
�r;�(<��g{�>s�����
f�\��kZ����nٶ<:�Vc�G
�� �d�֯P ��ӻcUX�7җ���I���v#40������L�
�e�\�IA�5��Z�i����@��Pߞ1M0��`eb��N���}�0����xD�`��}���_��t� �T����K-o=�F@�� ��gW~��+�+���1``�IG�?�g�n�(蘳,�D˯��cv
�!b5wE0����
w��n�r�:"`ϑ>(W݁��<WU�zF�Uf r]g����J���TO!O�����W�g���*�*^(聊�YKG ?9|a#�+9���K�J�aSԜ2,=)T�m�nx���p�<Ú�{�2�脇-Q�ly�0�/�[M
��,iCӆdC}B�y�����Mm	Mm�چ��@+�`Y�h�� i� 6��\��h��Ѡm�ܝ�M��:�^,��L����w�T��Ƙ� �ǋq2M��7�1Â l;�CP�-n�OK�J��i�
*l���9ɷ���볌��5(W�=���"�NyC�6a�9��4�<s�^7p�"7M���Y�3Y�UFM��R<HH -\�����4��冂aTz-WW9�QZߑM/������'���Ym���5�:?�����.Q�CT���Az�n4�m��D��1���²�s�ӐuYM*��7�3`ι��P�\-EE��t�E26�x{k(�B��/�s�6��kv� Wbh>��l�b=��H�G1YB4Oa=~�C��į��H�wZz*4rB����s�XҦr�խ�������쵳~Ŝ�1�:��|�-T���+�R05�'D���/i�k1M��2�ڔ:4��'\�gŴ60���<������o���($��|�U�����\���ʡ�O���>�JMy���#�Aj6GvOAu�R���N$����H����S��d�#[��&�9g�G0�*���Ej�I
�-G\c��@�Vp�y!��#�F����Q�`e���4`��/w2�E�����L>^xc�+{׉�;������n�_��uBQj���dƽ}�;.Ճ��c�T}W�n޺!�+�� �D�Os W�c��h)�`T��޽x�_���ė�ݼ ���{E��P{?l/���<����R\j��88\���f�>gDD��<���4�d@1Y��6�l�q��ൺ�N�e�b�a�6�p(��`�BYR�ae�A�����3�]��zļ�$�ѬY�2?���n�8%�u��У�/q��*!?�t�$_cH��l{4:a�j����&Hw%0������'(�K�3��Y�ڳN�����fY�����Q�:��O�r����n%[Q#.�=z#��ҢkSo�(��ɺ/2��ۣz@_ԁAS�4׹�;[kkojc֗�+ϦTbp�޲2�*-l$;�ٰ;P�_�/����n�����Qt�'�����;b����H���F�5@���$r�a:��$�{��� GF,�sh≟��{�R��O"�:jo33�Z���	^��	�����jJg�����^E@Io���
H9�lOEŘENJiBj9��5'����d9�	G��Q��lyo�Lm_�X�$����1ɍ�6{�O?M�!��M�MtҶ�X-͆B��ro� ݗ{S��߱���#`�H���6�W�i;�}P�י#���z�gD��SM�ba3�4�4�x�ĸz��..�����^}�1�U}���,�S�}�s+�;pDpr��$2�������(\=��)w�KR�I:r��e��A�gQL�V������Q�o�c��A	j"��#5H��l�d��r$ڱFv� C)�n4T�}�^(3��<��;곐������g�z7��@e+^?7�w��?t���Z�ۚ��D��X.�5"�Ů�c	���Ί��y�I��u'��7��?�_}#K��6:*6פ�R3P�}��*�N�9WenBY�/\��M䈼<�]nDL�?٤4�wM�E�lG����.,��2{D�7�M�Ar��R��� �(lГJØ�W�l:V�;-Q?u��M�ꟜID3��Zr�g��|B�Ű�~�Y�1���u�ӯ��~����3p+ �h�Ps��G-��s+Y_�z�~ǀ��R P"|K��m:x��Ž�tե��g�����<�Vw�:��4���=)Cצ�Ɵ�XL����`��̦��t��-��q`�%����7�k�`9~�k>U����}�Y���nj�zB�	Ⱥ ���j�G%�4��9�g��#"�.M��W[�%��jT,�Xj��Lo�)^H���b�
+��_t�M:(t$�Ѭ��XƘ���)/�)���Ʒu������1���'�t�\)�/����N�O�֑jW����rWi^�`��žb0���=�u!��!Q�T�%��&����+��\?"�C c�{@�0M��{z� ��=� �\��7��W�l���t�a�צ2l�!G�ݴy�K:a1L�[����� W�}�P^qG�r��ə�S���ZT�ds��]}��5��\KQʺ��>>Mn��o-�|�^⤯�nZuUi�rp4�g�~�,}�+���%�Ĵ��'�{�+�A]���<�8g3û�[,./%�7X����\�#�t�GV�%�/DlT?d�*;�[Sj�6���l2\�@`z!�^CSF͛���@h�+O��H��Ű�\��b*rw&�<'OA(�=H�^�{V���$����	���0��OT.� �[��K�	y.A5�Ԥx�L.)Z�V�?���/|�P�	�$E:�+�^��+H�t^51#���s" ���p��U����F�V`3�yHm֌#Ml��������"b,�#x�c�H�0�rI�^�}��L���=�K���67��lB`:�GC{2\"���+l��i�C �C{%�Nh&v	]b�Pg����_>����u�R�E��+�f����Sw�����C+]���~O�Z��0o�z�����[j'>��(��=��.I�g��`qT��X��U���t�U����$�	I�(>v����t��NU��uRx�K�TP�|u�d� T3��!l�νA�3r�v������d�Y��%�oL����˜XZ�7���v�'�= 	Xd��/��8Gx�cǟ@�=k��.!�}:����}���o#�q�-�*�ss���OJb@�;ju�M?�K!tYS�
��,zl���7�t��x䖼�' �n��9�Օ�!ΰ���#����J�K�7�� Al��F"�`�4`��k��`�����\~�y��m^K��<Ԣ���X@OR48t�}dҏ��M��°��Tl/�׋j��&j����(�,��>��y��k�ۧ=�pc+� �
*����0(�sD�QS	��Jp�⚚�H�RI��ν�h
�P�ְ�7��H�^t'ls,��ȍ\���{���{���;�c1��z,���R@��Ì�"����������o/���6ڢ���Wv�QG/��L�,'�
������Ү���K#ħRe����J���0)j�\���}��~���z�Ձ������.{���Լd����p�V�dqmW�G��V��e񾿘u<��"z�Ѯ]<o��-�y�ލ�`�~���f��ic��5,��~W�[5�����~�X��f�{����X�q�7�U"���1}�rӾ���VT	!@�1��l
Ч�E"+�6~��Ǣ�-k�3�&��`���)p��g�du-�Q2�9������S��}F��*/A�m�(pWIr
b9��i
�(pc�ӻ�R>Fɲ'��s�)�fV=~�/����0�M=������=��:�o9I��>�7���7�����~?�j���*0�g8���S�{������U">��a��ʫ4S.*��_IJku�N�Aɂؼ�xE�J����/�E��ٷ�fb�s�iW�z�U�x7�I�o��K�W|�������Ϯ�!��"-2�7_G�Xj7Gk��(�C0�w����X�� ����Q�xG�%H��N`��ڒ���ɠ��9V����E��u�,
0�d>����J�C:���^�Z�����+�.�E�q����[4�7?�1�5�����`��K�`]�m�/i��C����T�{&5�i4#�ݏzy],`�r�2۽ۻ6��i��=8H�G �����G�F̜�"r���/����5e\$x>�@�qI���h�S%�=p���#X��D������{|n%�7�/�Vҁ$i�����{��x�S#e\�uP$X@����`�������a)�D�rgȸ_K�UCk�Cq�ں��ͺ_Ud�����D���_v������!�4V7�\њ�5.:�9q~��X�(>���߅s��ޫ�4�c����G���p�ڹ7�Z8V��!�S%��\Q"���cԵ����+á�bA@GQɆ����
ٛ���02���z��o�g�|�
�оT�Q�R�4�.�b?�����m��p[�ﰹ곖ڨ\�ԕ�&-tL�Ҵ�F��&$ZZ�\ܺ�"LW�S�z�?K�{�����-u1�0�E��6�,��2k�jE�<FH�:=
l�B�6�W��J���B5txV4*�6���fϹHӅ}׼4��ge�٬~����c���k�PÌ������] ��8�-r��R>k��9�����>˓����8���߉R�[Ǚ���1�V��P�e����e��'P��*Ō�c��b�I�������oy���ڻ��V�3����K6�eh2��pD�~^���;�.���{���k	i��쁋� �~}pH�i�l��GF/}����eD/e'��ptv��bc��{�����4�E���K����(�p��+ ƝB�C5+͙o��h��p�vi�C ��M`��
�t��?3w4j#:�tY��;�,1��mq�,6C��<ވZr��J:9:�+J9��E�P�F�L�
J�)?z�c[�嵿A�+�*��#�#0�Z�J$
��9�Un�RhS�p׻�I����m���T������C*�)��x������D��o�!C���o�ލ���xW-O�`FmKn���2^��bіu`�}F��ӈ˨+٪��8����=�H�qVZ�u�'mc�vO`�
�o�'F�v侦ŏ��$!�C��י���
��,���6Y��p�i;X����!���.;ח�"��{��V����,�k�'of��`V�$��Fƥ�A�+�,��r�̦�a�S2�y�^��B`�s-�.K�����a.SOk�iũ�Ѹ���?�q{���mx���b�n��UQ���+[�sq�nL][�0�@{�j���6��X�����_;�����p8�p�F�*���N�JQ�{�{��犾q@�����lRSS|7��"d�D�P�����fX�:`�
$z�u�wj��TXc�AL�D�A���$ơ��'��H�#N�"����r��X|k��#n6���,4��v�Hʳf�5T����|�d�W�M}`����6���jq	)�|�IS#�P��� �P��<)T*ȱ�=�Q�_��r��@چcȆ%�=Y�T�����p��Tև�c!fFi<P�&1��Us[�%���	�T��^縗Xa�9�k'e�(헆6bEڣ�s׏ 9�f�Gv�w6'^��5�����t�Z-�n����:��:��9r���*P�czdK� +��D�8��䪶�a��S|�cs!,��5��Զ0�`Cux.�O4��3�:�t��\Ο��;ŇH�$�tg&�08D5Z�,;��e����D\�1VK?t+�%Ɨ�"VS.m5P����z]�xLy�PW�p;=#���[�g�ךZB��Т\�qGz7	�iv��E���A���q��u��j� T���v�3��2�cDy!Hp[�td�>�s
�
@͍�M��O�Cj��7�e�ח>��w �w@E����8xz��;3e�t%�?��F�#<�P��{�㔓f�������w����!�d�<?_��Yy�ti�+�=,I%��l�T�2�k��wS�)��Ќ�Q�X�:�{��DGm��G�w|�4֯���+�g�[S��n>(�1�9�����2�Q}&�����-�%�Z�7�YO_�sQC����8�]E��=�	���KV�ͦ�{���&l�28���V�fr��5"t�/=o�.�TK!���rr*Z_ڿ�z��H�,Y����:�C�\ߍ��+�S�X.~�\%G,,���@<�aL��MR
�VT�|0H|͸�(`#����b} �T�QZ%� �[@S[�/Q�lc��?)���7��U�-�cN�>���zK�i���
�A�0�x�:g׶���Ǩ���Z�NK���6����2D�}2��&i��1��`dp�4S�ɹ=R��J�C��{�G�_�v���/��q}�^jL]�z��*[fwW�0K	�]�4�f!)�g���+\�C>V+x�ia�dt�u1�a2Y~��+�;�W��ёc��'��Hg�|�X��9,�i�fF~F��r�����/���9��t��=/��BV ��zc��{��˕(3Kq���Z;��J�e�4�0�K���6E}�j��G�	����6c�ixqJ�^����gQ8����rn9Z�D�+��	�kh�YF�G�y�l��D�PqD����2o��J���,��;	�IW�dԋV��^Z4gnq�"=S��Ƌ>$#.c��vwY|Z��5����y�!��c�
(Fa1��m�}4�\�Ѧ~�p�jڗ_#p�2�쉒������9���@є��:H%{���c�a*��g�� �Mn���4N��k����3hq�^�ox`��i��i~�B������O���/OmCֿGER��&Q��BTӁJDn���{��C�ZgaE�XH=1��L>�P��1uXB_�^�3yy�Y��������p�(��N�t�����}{t����`�`$S�
��'��B~�JO��T:F�p��E�S�pr��(�(�-o'm����k�t����X�'GK�~6��%�'b�/�	M��?��{��9|�9�3��	��	8<���}"�8}b����/���.�*;�/^�)ѴN����~I��'����ܽ,%���kt�㙪�%�"a��4��J��̎uc��:�}���h��V#�{�}�i�ߵ{m�p��^ޘ���!I�%����ٶ�PH�K-���'��d�l%3�8!{�l�7ޥ�X>�Z�U�����r��})E#=o!�c�-i��1���z_��n 9/����n.����;�y�>��kvp����%�bӎ�
+P>�.��m���wD�61�7KKH�t$q�ª�9h�s�Ԯ��i��Xڌc�v���22ڒ~�&�֏�F����D��Y��W�TA(�u��z.�^�7��������g(*Pތ��%�v�����L/�|�����X�������`�R�%�`>$	�^�-��X^�@�ɮ&
�l"yi�*X�a�Jb��!G�5`2�I�v�c��Z��e�㐍-`x���g�n����:'[{��� �"d�,{�ù�����X���pH�h"�5MڰY=��Ѿ�Uq�Gs$!�t��s6B��f������hiBtu�wb�ј�L{0�i����G�Ce
ٖ�b��+���8����ߕ��p���Ǟ���uN3ۈ�C�
^P�k��_�f]��꧄�Ԁ����ܨ�O_��q,��ܯJ��^��z�P�@�#I��*��!ߐg?�a��\����{�<::⿝�fZ�̚r�ϸ�Gh&��:Ҿ�K[��47��E�ղ�G	r��Mn�Z%���ʼR��R镴	ɛ��v��ZC�ʫ�c�;��;0����� �Z��?[�3T� {Ĳ���J�"fϸ�7��t�lJ��J�z����j�P ��0}�M."�G�B��l�.��>��Oom�5�_)ؕ��q��;�y�j��i��Q�5ZatBF@Y�%z��?��ݷUkH�����O�d*����1���!����>4�Q�� �l�+PE�~��2���jr�\?q��x?���LH��>�iM���(#L����=z}9`� V�BY
�3C����ӱ��M~Q<FcIv:;2� ��)p�96g�A�G��7�x�Ac+���띓W\Ƭs�+ �30:���z�Z� Z������+S���?C�@��oB]�Gט�����Wn�ɢi"�����4T�b���ٶ8���4u/'3�����A�R�8�b�B�;$r��O2�ml�yF���!�����Chq:��k�u��/��<�x�w
��|�:���o[�G`=c�W��2�����{LRpT�h�T1?{?X�Zi�^�څ��_������/҆p��-mX�G�\�I!/�v=5��edݏ�>B��/��7���s���5'&��ɰ��R�[t�!�>ԓB-:8�Y�M��k�D�}�(��
C䟜�h ��+���cp���o�7�R`a>7#jN׉���ˇ�F�>�g>�:/?i3oq�Tw�d��A�sc�6�Z
F3��{�=b�a�q��M�+?!��p3���*������/�E�7)�Џ�/r�r�#��@��)��נ�b��I��x��/K�]�cf�X5�����mn��\@=(
�W��-��K�C]řb��ǀA?��q�z'n������LfSs�r�%seܥd�3�=�l���dpm�(���J�N��J&N�� ����S�KGȖ�{ ~���:�5�nz�'��<3R�%\~���L�Z2���A='%��>�v�;���C�ۯ.�+F�ծm�k�)���0��_&��I�|��G%b����ǌo�r��e�o2����G����v�"�J���������>/��и��o%�Kꍐ��%�i�M*���l��E�7n0�uw�2w��S���jo��Bem���4�m�?�`�ْ�q����V�A�T#���s�6,��B9�{V��r�N�*4/< ��v;QB��,"&�jW@Ü�����yXA��%^6�NE��w����X_�P����Z:�ۺ.���^��v��}s+l��+��J���r�*(��f�����'�Ϸ\��PE�4��iY�O�8H�M��j
�X,�t�%=�
����z2@��_�M)"#6��C\ ޑ������W�?7|T������j0֝�{��P�d�GNJ��H�#��	����aO z��~���[>B;�^����K�(�`�c��5��4)\��rkx,��X���a��gWF�����foI�e�?�,��a�Sid�{��T�T9�;�0*��a�y)����9&	>��G(������:v�e�t9�=O�.��$A��~������p2P+� R��ed�k�܀R�Y
���N���7�P4*As�K9Xà.Б&Y>�l�-�$|ѺC��1����٤6s_5t�%}=����>�[1��ܽ�){XKP����3��={�%²#h!]dM�����n��vR�TMև*7`����<�g�f�391����"�����G��PE�/�.�_g��N��1H�cq9��5L�ư�!k���$-&��[%a64ԩRY�K�04�!q��@��d�9t]Ы�f���wwq�a+��4�uA˕����{/�uF���Oo7'�:�ve�8ڃ�ܿ�Wy[m�4M�s�#Z��_�
���^T��&�2w� 3�7���p����Q�a�v3{a���\���F�!���"_�� {�_�^���!]���sm�&������hʲ��N���K��I���,�t _��(b�W]*��Go���Z&F�J튄݇�'+���M����@���%��_@��y8�*YL6�9�݄��r�(�T��2r�����w�	OAL�[����hYC�`Gn�����1�$/��u�#��d��^ђaECa:J?~��X��ӿβjS�q��7�+�-��N�ob��W�k�K��iS����8�UN���|���D�D`���i��?Ks��$�c����wy�S�����o�8D�{��h%�Q�EK�D})���.��ʙ�U�s%�L
!-%��ע#�'�?4�
�qP)^b@��~�|&�V]����?r��\.��BȌ͘d���.��Yi�CT(B6�,�����S��g����ð��|Z�zSi��V�����w�$Y1H@F0�^d���Wˎ�Y��Aa�/��)u�_}O6��y�d�Q��8O4a���7[�<��O���2E�=l�B|�ɧ�~f�B2�ʺ��� R�="ΐI�&�o�!\�}[Z/�_�Ju+�0Nťh�'�L�V_ RM����L"��8)V[���uK�߄2B?`K��G>��L%݀���M]��=n;�N�̥RU���?4�x�YH�KB���E�^��/�H����
��t�\Pφ��<�.!�#����^����i't�#�/i\�r̵��P�l�Tua`5�D=W+JV/Q&�ⅣU>����_�.n��q���4�1xfо�aڼ�K���}p;��]&�ɗ싚U�A�?����!�T�q؞B�X�(�O4�=c��=3�8m>Q���d�4Y��}�Ք&K��ѐ�C��ڴ��l�L���S<�����f�㔶��;%]�^Ow*~-N��1�<7IRkI��'�Y��<_���]��u�>z��hkD���`��2Q�q�F�tNF���5*k؊�M� 9��e�5�R.���U�f��bͣ��8Ȃ�n��x"Ս�y��#�=�"�yh2in�cY�h9�$I��
)�oa�Y�\&�t۟��qd�z�e	T{8��P(G��Ũ(֒���(�Q��Wa���)��/��ɐ��_(k��W���a P�l��G6�O��VR�ǅ�M�m��~�7�ɒk���\�,��A����)�9	bl�.J�N�#`�/?z)�� ����i3���L�r?Bsp������ ����u@��ꉗ����#��!5�+�y(̄�W��*6�G"���o�V!����J?�t��<=��sX]�G?�V��6�"qEC9�de#zo���Fm��S�^�ߔ�S�@�>��I�V�$.H������jyx����-r<hGH7�~�9HkBE��@t>�H��ǆM�3�P(��۟�~n>x��z���4y$��`E���p��o��GZe�H"-�C��nt�����ѐ��-� ӟ�T�a"�fD���׫�J�[ɏ�������h��b��l���F�ihI�Â��l�v������'�l/��X��7)I�l�Y�7�7�p���w�_��o����/��������Z%B���4#~󊙫�(6&�򙾡iw��u8h�R�S��[���.����JX|~t-��qvd��������=a"��!��f���fY�A�,"*��~�RGl�9FMy��e�҂��%��a@7ۺr��$�qDi�rv���������Co�;~}�D�A���� 3�3�bd�'f�K,[��h�~K�]Us���)��������N؎0��B�9�ő���b+���5`����Y�D0l~��6!�"�4a��|]�x�fm5uS�k��!�7�Q�DD�M��N/W,uܹT�_�Ք�̧K�-vtip�ŕ|%��� P?��ӺÿX�����9q"�7�h)3�KGD�k��91��ݫtM`j7n-;���} ���aZ��h�D�*���=;�t`�)i��J����8�.s�t�Z���Lȷ��U;�.6������a|�+c~��"�y� �,d��?��ܻj�I����N#4�-�y����C�Rz�;R��T��kf���^F�'�^ ��NF@�`�д@-��ʥ~��������CN,Q����X����M��~�c�$ʶ{���a6ʫ�θ=���L����oǳ� W1;$�\<k��0�ru����>�tJ�ᓡ��E?ݝh���)�ֲM9�j??��k��]t1t�:�,���l��
`����H��2>���;�X�!L.�[�"4�O���X5�Ի���T�^H5v���.F�C��١g�#cg��Mp�6E�d��\9@�a�}��ZGD8�*V&�	y���\sv���&is�I�Ҋ&pG���6xF�$[��.фodU�]5k�Sr��7�t���>IrOv�Eˆ�F�߳�Xs��� -���&�?��m����5�QЄ���H�pn���@�C��[�E/�G�W5�+� ����j���G�{?UM*����P �9���4��'ن/�!��;�آx*&��'���"'
��0�v�S{���K��0���f�4U�0�T�	,i��I�l^��u��~�!M j�v��h�T�m��h�"E`V*�}s����B�Â�E����Z�CC���R��8�M�[���8�ME��	��ʸoVQC��5�>ۙ�D�Q���,I�>� =
]���K�۞=���e:ȣ/D�v�L�R�$�ɺ��l
����I�ϭz��⡹�	O&$�+[k�c��x�b!9��E�^2;�ި�y`�����Ȭ>j��:g�@*B�������_	'�����F�O/n�[	�4�����tj/}������ޞ�4��
p����6�� H�T!CA!���-��/to��M��ֹfڰC���������q෡�ê<��B���� '���X$Z�X�+B���+7/W�k��hf���?�?l	����u�]��\��t֝.m��z܂.�ؕ�j�.��ʍM��U=)�i�̅�@�b�t��v4�!k�w]U�г�Ȼo>�[�����Kh��D&_�s?�l����x���|S넑 �y�&�.^aF����	��Ψ E6���B�_�6?�ui��V��!k��d8l��ϯd��t�.���\WM�}�j�:���H�!���D�5gБ��=�T'��W��� pC>�~j1����E�������]����e߈��<=^Jtc����	����<[��.g��;`�����q�����K�>?�)�F� U Ad9#��iG�w��|\3��Ξ%ĐiC����QJM����n�,e<TپO���g�q~Gv)m�����p=����|���Wc��yA{@@�������������>eퟑ��x0�0w~k���b�y *���^�ݡ��Vxr�X<�H��.~����N���"�dE\&�L�kr���|R�P �я��E�K�;��7j��1%�6ݒ��yH���l��	<�yW��t-B]|f����OJ�i}��z1!?$����!�AE��������C6R��U���=�;RP`��>��	��n+D8	�������S�gw�@��<eWk��Y��pg`�ҽp�cQOQ�2�Ϸ�_��A��{,/����P/�jY �P*��?N�MQ=��!:�xEi�3�^�g��~�z�I[�@�S��G��K�]9�ҏ
ŝ��ֺ��fpg��P��M!�3K��,�)��mU����鬜� N�s��m�d�͞��J1x�:�9�=��\�ѶH,����$���JI�����W�d�NCSU�^�3�l%��o�C&��Q̜�{.[%�(Z�,����?LY��qy��.P�L��SSE��u���je~�F4P�q��(�n5Ѽ	�7Ӳ�͸u��,��co���c5��%g�����prh��N#���I�Z��@R��`Ĭ�&#�q�+�0�^�X����3TU�	�l�2l��d�5�"|E"�6�F��T�nQJu!�;>4@�e|u�����p�ko'b��o�����P$�:~\[���M`b��B�:Re�K���^� �m=�����5�n�w|���!9�I"ؔ��c�������F�Me�	ص������%ށ�fj���w#e�¢�T�8�zIy꓉��<|�#0�Κ�!�Ufx3���[	�"+ ��tB<�)����+R�_�uRѥ��(Xg��@�nb37�f] ���������p DP��̂P��gs��N7����3�$�t����x�V�����<���u�
�����d݋�Kj!$+r�Y}�D�R��ݻ���_*��i:Q�G��Y��:�K�����(���эo�U�<�
��� 3���i9����)��2��x*Dj6N �uS��~0�U�t�ԡ��+3`�D� m��,�ex��fŚ�tU�,N�5�p�!)�cQ@������M�ӟΙ����B��ިȢ��/�T3>c�3Ƕ��ş%�JG�%�f �y����\u�P�DZ������PD�ľ��9��(��!�۷B+<�?c��{��͗z���-�tz�F��V��A�"�l�L����UM��
�7k���(y���Ib]�������Ξ3���7;�;3_+���6qL��L��]��/�'�<��y�{�^��8"�d�r�:o����g ��[U�����J��3��ۿL�sT���L7��~I�)���M����k�G�J�}�_��`�{QJ��<�0c(4���@�EU��c�b+���c�@���Hؽ$E��&'����jkd��U�����z����y��R	�>�2L���۱�آbRƢ�چ�ŭ�����|Vh⿏��
����m�]'�:�����k�4HWOS��$�Ź�:��#�m>��]�O��c�����T��� �MUk�* |H���K]�����@��Ś��Z�oƈ�+�<{=Fq)���,GT"����)G����)��*���`@`�tՁ�m2-��V��w�=:p�B��w�ªi� D���r�%Ry��c+HB�!S��{���V�P�w�%&Bu�a^"��.�h��|�������Rے���{��N��<�=��呵��7�O�b�oH�s��.�b�{�����7B�AD޶l"�L^ ;<�z�z"��H��{R��?��v~���=cx�^E���6x�ux$�:�ҹ�$%f4�)p���v�Gm8U�Ձ0�*J����/hJ�KT֊�L�7P���F��R�jҦ�M	����G	U��^���E�͢�'�ߖ�3�/΀I�˓VvAls�e�$r�f�A7E,��g�r@�h/3J�ީ���� �h~nFF��ۘ�H�2�"���:�`m����T=��0\ycښ�B�NӚ�M��&{kl&8�]��ޘL�@'Օ}*x?�����v+u-�&S�u�?��9�Xg��d5�f���͘(@�IQ��6��J����AD�3Dxe0��-��u����5��`�n2��W]e
o��Y��SG������`�
 ㌴�M�3�"�¡Y �A,s�$B�ЊG�&�>�3S=Ng^�]D����)�h�%�\�׮A����9�`�V�b�ηɢ8��\F%���G�u�����/��M��i�+�Ź�/����5mZt�1�_YQT"��=%�M��$O>�w��#�t������ᠸ9�����{� v�N��V M���!��bf�&Kjj��-�SE���v����x`�K��To�|!(��ʶ�[�D[���ݬ���t��0�������~�g~sI�F��6�`���2*F�I�X�[�3xU�ʊ���.������F�q|���H���v��2�4�F���Ĝ���7gQ�4�R��z�e���|�,�`+T�ב�!V,�]�܈W����艱(�|tt�����]�)�E�>�)37d��R*3M�y�C��+Еc�5�
����G*��B��t�1Q/��lI*Je����	h��ߓ�I8��G��_�M�RV��������_D��f��'{
�)��@�\o�ޠ��?�8�C��W��C�Q��p��}�U%�o�]�+tt+K��-�T�C�5�=�L�f�<ħ�0a%Y�S�0�!Ff_|l&��}�����9՗[HVӎi�d����3�홱Q�<�X�<� ��V�
����!	�B����(*�	�	��Q	�������2�A��:6Q�"��x�0m_���٠o9��ؖhm��q��Z��K�x�3�¿�ͩ���l<��k`�Dl�s;8�(7D�nL[�f\��b�:�o����Wh���p��FK�$��F?"�473��#
R-6l���A�)Ds��Dp���E������?;�u���B�#�¿�a5z$u �~�;���>���D?���H�w�������U��|B$h�@��u�[�#�9@9C��;%��~�}Z��0;/�̮�����c��K�N�D��u��6A�E;���g?Rl�<�|�� Mb@&�Ey��$�^'�/�����ݒx߯ d'���\"0�#���8e��Msm���"^�o9MlQ�NjXJ�����ײz`������Aԏǚ��S��f��b�P���e+j���G�w&=����@⢥���7�A��щ�B�h>����g�_�T?Ӝ~�fO�"���0�x��&�B�R�G��|;�j8(�iL#�~3g" }@2
)���?3~
���+		��y��r��r���`m'����J��C�|��������?Q�*a'|���l��������ov3P�&�-Ef��)_��{xQ���+Y�y"��kl�ǇV�d66��F��e�sR+�|�ܴ(�b��^��I������1^U��ɦe�Yr�\��(.��-�62L&M�z,�6�W@���y�2:֭&9�d2I�φ��{�g+��KV�,�/b��Sz�]wc׌a�f��g�XCM`���O2NC�����]��7�{gl�^27�`uV����aD�7]}j�C��d�WEc}>p<�JB�x�iXR"���b�W'I�:��8����,{��F�(9��b��^;���8���0g��o��H���V������f���Ȑ^�^�k(��� �&�X�D"6ר��H �
t��d{�ڹP�`?��?�k2��y'ʑ�M~!_9���8���I&d�.�
hR�����"�0�Oj��/���_��������c]��̧�ָk���lA���	��Ax+�7��pO�����+�Sd--��i��a�P��A8����&z�am��r�),yoԮ�c��(�*+��4�U���W���';g���)އd��6.��G�����@k�Q�r�e�Jˑ}�*>��f����\��.[�KH ��wB����7�	\�����q�J�qn>�b���2��C;j��kⓞ9���C����&M�D�Ma/�jWگG�a$�����[B�K�>#��kw���gwҰt8��𲰛:3SMVyB�"�I��Z�ٰ�H��|[B�
�.هA}��XR>�W����;#�lӌK]Ě�W�|�� L��L��3��u����Ed�i�����1�Ӗ, ��Af��Q^#����^��pj���[�2�����QZ�j��H��m�� �@�K��{f��Q�2�h��Rj�A��5V�N(��V���¿}�{�'���_��ʕ���QF�=�������^�W�:�op8��ah���j�>����GĤ� �`V`O�L?��'��̖�U�mj��-��?�$B���n��]����m�υ�%+<Bl������EX�ar0�x@������"\�vbH������r���nw)S�����!�ϴ��J����z�:�O8��o��ڜ�eY\����v�~��V/fd�ZY��6���T�ߞ����ai%�fLk�%V��GQp������T�݇�:���"F������^7G��m�;b(�d��5���D 15�����^����3�v��=j�1���u��{�~�/2b��Lӻ����R�:�4�W�s ��%�'�4���>SsH|d6F5-�#A��V[ǘ��w=7��C�o�T����Q�{lsAk�����X۸�S�Z-lg���"U1F��0g���������Na7������,fN�Ü
Iٻ�/LJHa�S��p�e]>���WOE�A�j��%���g��?��E#8�Dg�6{J�TɕY�tWO&Ɇ�2���.c��p�ʑ,K���؟�Ub~3�ڃ�i!W����қ%>1�+�ȴ��!����[Ml��2� ������E��	y�`�M:�}0g$�[���m/��s����'��B�tZ�ӈ�u�]b����t����z�z-ʴ��V�+��AC����� -��#/(x�Ɲ�n�7�qG�u��pRw�����9��I��-�㖝pj�*��7��W��%�I��7�&�N7���b��x���M�o��;��p�Z��m�]��Dbׁ��U�˙N�+�B���>�s�J��J�΢�<?��A���7���c��8�6`�d��� cVC�~0���.�ڷAlv�j��K���eOn��������׼�����@��"Ȃ ��VT-��y���@��0s�5ߖ:�����������t�Pp|
xcP9�x�>|���g�<���Om6<c��2�Q����Z�1�R��rSl4���s�Ӕ�܆3p��,bk�Ѫ���?�]�����I�Bה�����)����*;�."���KBM�N�g�jyP,x�H�yGuW=��(VMJa@���	��6�C�5�-���I���>oŕ�E�$��d�A,TA�N����~'~X��t���dN�q��~K��1Ў�Lv�dQ�ix�º)�Tme�|zK�@o�f�=�ʭ��Ő03�Ӣ�� 7'iZj�D��=�UVe�R�����{� �-s�]~�ޘ�ǟ��(��
��&T������/:
* ��� 9���vKB�3�s�6"�쇸�6z�~fܓ���Dju�0�Xw	�߈�z�>�Y�����y�搫��?�֙�>~ş��8� �^+�o�,��c�܁\7���m�LT�n�JdN~���ѴF��K�����c�WG�A��d�Ja�n����?�e#��t[�?R����
�Ǌ��-nV\m��?�/�p�s���[�K�T���Ծ�C� ��A7*S� +�F���U_��+h'|���"'�b�i����4k���jQ�
T��V|�b���iL�1sp��r�������B;���sRb�A�_L�����R�JUzt�[���jM���B��<,�)��!D*����}�� ��n��=�?:��ͅ�'/�d�o�}��v��I+Q�ӂ���D�!����l�jI%9�Ϲ5��2�ſT�!$*1��&�Ч�˰�&�Do����sb��5��{�N���9eX_^Y1��N��WSf����;$�2ϘM�;T�@$�	9��>d�$����]lv�)=��c��.�M]q�(����n��Q摩N�y�p<rx�?��2��n��׼bsJy�����5�/v�ZL����;if(�巨��4���w�4e.�}��)�Wo�r��3P�f����E���7%\��l 2(%�2a���=�V�6a����ݜ��m��<
�V����CB%u���Y�cVP�(]>�,�[d�
^��έ�]��</ت��
�/Pˆ�p� GY[T���ܸa`�K)��8W��e*��)��h�b�nz�:w�?����>�!�.oϝ�+��#;�1%�9�	S�L���נ�Z=�Rz���{� �K;���	�����{�i���ӺT�]1	�ixw�iW�D��N�ЬqӁ�7�b��f�[ڗ����lK�o���S����ٿ��Z�g|���l��������/�j"�0WO1a-҆�����#Y
M��C��R������?I�VAS(k�)D#����ۢj��c�k�W��:]��G�_�?���D�;�?ji�@<bZ�i>�3 ���{���!s}�1�gs��m���Lۋ��W�Y�2̂���D�p�{#%X/M�-�$ǻkQ�-�/������xD}�\8�O���X�U���:�SI���6`�eadA×���i�9��jYL.c�������&��p��i���уNʎ7tV��?����e1i��a�:p�J(�:����]xÜ���<�o�9��i�"l=>ƹ4jy��&�����F�����
������L �-\�b�)�|�js�B$��=���D�,i.'Or� ��e��W�C��3���d\=�+�� 8�2��6��O"�,$ ֕�ݳZ[BO���u�EA�b}����=;BU	�@q�V�ŉ��y�ѱ�+A��'��,��;=� Z�j���`�Bvv]hUݜ��kn��i?+Pĥ�?+-N�c��	��K�q�Gf�`�RO������DX�&��7g~:2�zl+�#Jt�Z9���)'�֙Qi�s��'�V���F
�o�s���!T;�L��Q���Hx�TB?�{��+zSe����E��82�X�S�"{p��/5w����>������3�
����� �-����������㾦�F^�1~+~�_�D�ڢC��b���FNs�#�_����XA��
������i�ZAx8�wN�dD�N�L��6��z=��,���%���%���aX1R�7�^�]�����Z�n���:Q"뾶�:��L����x�I���I���~4�(m�������k�;�FdH�i�s������^��85-حd��xBPNî�Ƶ���{���|M���H��#?g��E�6>9 �D�Q� no������śR��$Tψ�j���r+z74.��9����P�d+��V���Si��|w&zH�� 4C��yx�Ɔ���\�N��$��`BGl4R�s�Iiv.t!�w�D��N~r��é{�uM7��j��l�8f៕H�1d���j8�Iк����d��/��YO����[$%�n�_�u^�A�����߭�����;����l�\�=qMP�zƏ�J�i'fh"I�s��s8W�����H;�3�X�dL�;1��,1
� ��Z4�[س�Jn��|��S��CL=������ǺpDۜ�a�f'���J��
/��#�ұ��;7��W�q��
���,���݈��!�{E��@j)y>J�Gk�~@!�ؔ�y"Y���g�-�Ɛ���0�vG���,�_,,��D{W��m�y����DㆅݹW�������@�[��b(��鿋��ԽKk,�vVێ~�/e�>�9�]�QWO���r��ߴ�!��ɽ��6��.Lq�xd��N�dR�(�9�_�@�8�Z�/�:2*	n&��t$��c#`��"��ލ��!�ɾ	]�wH�h��f�Ԝ�X-?�p��ᙙ�#�&q�PY..��%���Dt����,����C`�s�"��iEo�KDDZ����+89����d��{[sz����R�b@*�Ƞ�8Bj �*2|~6O�J���^^��l��Y_'�=4���t�1p$�t�݀������T-��z�E�
֔e�^ w�3B�8I���rrG��0Bm#�ZI���ڶG�����3��cV�N_8�ŻX8���"�����,�_����A��U��؊���������?�"�F��w埫Qf"�C���7Z� )KO�æXO<����k9�(����Ś�� �q2t|�h���5��$:������e.��
��G;E�Lf�pPx
��;jZ)�=��yNe�l���?}�`p��W������T��Zb�]C����8-��{=V�h���(鸈 �����)�T�(K8+�`?��K���f���p,}���;x���U���e� <����V���`FT����_?Rs��'��TS~�$LȻ,��|\��*Wk�2�Y�p%g�u���y�n?	 b�ڱ�`�Urm庠���m)F��w�|��NDS6�^�h	1Oȯ�G4�;%�WG�l�_�Xꮙv2�� V�&���L���F
����k`�.�*AeN�)���S*��R0q-��S����7���$��H����\����hTw�(�Nh]t����q�~(����{� ���eN����?B���@E����-�y���-�e%���D� ��W�@�
��|M�lY8���Z%��X�N� �}�"�5�m�KfZʞ]�v�&1����������T7\�G��i���C����q�*�}0���ѻ�5w�y����G[�Щ�^���ϱ�ޝ#����ف�Q/eD�p�ȼ��<Uz��a�M&2\ƛȋ�w��	������ZO����9J(]�� Y/����7i�"ڲ&�T�5������7�Ŏ$���_�.����WJ�P`����+���x��� ������t1g����'g0�K#�i�"�����#N��kq�AT=iA��KV=/G��u���Sn���by�Sw�,����f��ߡ�>H�tT|v DM��J�w��)�J*��M���b��p�L�t�P$�s����v7%Z~~ٷz�"�Q��_��D�3�5'o��-����;�C��7�_��*�C�7��fr�?a�vx+r���~
��ˡ9��������)�(<(�n�t$�(!�G�N�6������X0��0.~0V��;�j�M��b@5�h���A�p�cI��]3��V�|!�c�i���*F�L��)�7���P��ULwJ�y����Sla�e3����$���m<j�����<3�5��2�j���'g����t��z
o�s���{��TME=*�K��?5&�8'T�N�=`��q�U��������-�o�m�A�0��8��/jS�?M��J�3+�e���V�=���s���'M�;P�W���>��� �O��e�KY��Lh�ò�~��V<�R�K%��l��5���G�����˺��W��wa9~��e��F0�hpf�˽�A��WGGg��28�7�F9V�A~Pkס��F�E�	erj(�>2��+��&��xi7"y29�O�H�U~��}|�NĊ(s������[�G�݉%Q��u����B
��<���Q��2XM��ۃp$�dg��Q|G�	Þ�*ܲVe�謊c�̎��>"�kd����!�zrð�{
��1k���c!>��$-��Vgr�4a�F�u�+��i1xK	�|&<�&�v����Cմ�m�x�v�����Q����뷺/��
Tq��$a�|�E�G���Rʉ0����F�/|k<y_�Tj:��{�O�i��b�܁�S��}���[��L@TT�:�g�-gan�� P�$�%��@�-�S+:��:u.�ZႮ}��|@;�'~iN"d�� kK�u��Bm�r�5cvщC�;l�&��E�I�e'����r>=���.��*{�]�;��)��Y�q9O���g͐қ�&�)���Z��n�^C�֟f{��\$��ݴ�t!�8ga��^vJh2;u��O�%����d�$�vbP^���5i�.���W[	 ��x�&��[S�~88���~�����&��z�Ya��]I\m�}M2S+s�% ��@D~m{j�MK|\2��ReT��j��ֵ����b�~M��5����\wM.T� �A"��"v6|;�k��F�ܘ�I��#�ݓ��U�p��Д�ɷ�v��\Y���� ��Q���<�&z�J�>�0�qt�I��
��@�Ǔ3�\���q���z��5�[���Qÿ�����&i�"�p�fۣ�q�gfEY���ݿev��Yi�a��r&����G$!	�.ɹ{��k��o�g��|�p����ۺ*Л�լR�7��~<W��/�dCM9�$}�Չ��%�1�{u�{�SB�W�w��Y�"Kǔ�����b-P�×k��	c�c�b��k���KȪE�4́.�M���r�ז���'�a���`���@�k괫0��'���'�^{�O<|�C_�ˑ��sD�����x�j�q���ܟ$�͸3���R55]�Ź�3sP����Ӧ�X��dGj;¸Yf��
��=��o(�عu@���ٚ��&e6H=�1؇���R����:T2�:�*���$-���N��3jm��ސ�qx}#�jrn��+���ڹ�${���T̊3�����;��ѹ�����T0W"���p�W�����Ź�.�W�f+SZ4�O]����s~a[�.�0l2�7��;${d��?|)�q���,`.F� 2��e�T@{3�Ċ,&�|�]|�x��G~�eb;��]}��R�\;I��#H��L�	��>��3+>�5r���?�z�O��lbq����(�^
�S	�m���Y���r���cf�%�ϰ�����������X�����0�#�#fx�=,0pc��X�����ȼ^j��󕱊A%���]S��moώ�z���l���v��S��I��c�=zN�x�2�xd�~�B��w�
sY���(�3�ޘ���u��V��:���ͯ��=p�㯇������IO��| ��~RN��v�صF�3�m<�e��P�(��R|z*_{5vN�lp�	)��UH
R���cA��+�d�8�������-P\�$Uv��ʧ�HT��c�Ŧ�D5���'*��Vu؞qc�_U��ڷ[��ʒ�@��W�e�?�0�ޥ2H��	��E�:�K��%��;�R�rA'i�8�){�R��'d��&��L������:0ޏ
�J��Z������x57��";�(��|.(�%��	�4��[�t�}���6��jz��S�?	�7�[X~Q��7�f�l�W�[`I��ޜ �DL��ZA2"�\�@��?�Tk�%���1��'J���4ʄ��b܅�%7�$uF����#�̤����_h�.bŌ� �ӱ�.���R����t����)Vw�ź��D�U���d��'��0��]�{O��o�~2R/,]���i4c�Y0X�m�h�!
��:��;��%�A"B�, ��f�@ٷ-O��u��(�Eޙ�?���Z�]�4!���g;Y\��=��Aﵫ����^jN�߰A��Q�rlo��C���(�u��pkh
GJ2��40d�C֜[bN�ps}���G�\�t�y?@�69??�`�/t#B����Vd�l�(Nx�c$��e�h�LT۫Q���@��tq|��6>���<:��)�����<Ps�Vb��M#\p�`�G�.Ul�/ě1��2�ƸԨ�
D�8���9�gS�q`��?�G�FC޿L=d#=�Ԣ���oo�B�5"�#˹77R�z��si-*�@�����s�8�K
M�rh��([�\"���5�{�0>�yJ5Uq�c� �}Q����i�5��1?3��hC^b�L�k�6�	9��`)�˹Sس�o�-"M������TK[K	֟�~�pRԂ��*�ۧX��L�5Wy��ϋ�u���Y�.�8��N9b\i9(M�8���G6n�Y�J��q��"p1��[��EE��f�����cVē(}�7D#�Jh:���"�˃m	�h�w{TJ:a� �NzC_�eHI��2����ћ��<��)MXn�D{�e���M���?y�'����ϑu���}���ϭ�Ǣ��O�-D���-e�ѳ��7�!���*�~w^�����~��5��^�{<����	�>�졭Kθt���
:W���l���*7�.�
���^��~t`m��W1�"(�����XU0,�t��歯#���j��%��DCҨw����Z��0����6+�i�H���g�Q'b���Bp�(D���]쓯����[�]E�7?�y˸��N�J4�ѱ0z���������߅%h��x�
�t���Eb�4������b)��̕;t�k����J�)v�R����򃩒��'|U��Y�m�?��l/Z˱�]փM�W��W�ԅC�`7�[K������/������S]�`�~�`x�b��`]�z�6�q�29����\�)�C�m���x��5�zuC��o�Sx�E�:�譆#!�Q��z��J�n�K��)8�PB!~��ч�ձ�{+&U�<l��}8v���拞�?�q�+�Ŝ�;�9	���:Ub/�؎��l�ciN��G9#���#f����U���|p:��b�7�TV�&}��|D	�k�W'I�[8�`�D�aӿ�����zk{+����|5��
U�)y#�9�؊h�;�d+�X���7���Na�.�Y*�� �x4�0�~>�E�6b���ao�x~��y2@W���J�x����jU�6sa@Dr����*�#�v��\��|2����cϠN���U;ډ�9���dҞ�V��X��hk��
�"rU:��xqnU�ȴ������-`�q�n�v�f�Zn$�_���e�Gep�$�4��*C��
�
S�L�8��ۮ~�՞8^��(@�M���PUla�y�oDZ���(]s��hA3��7U���h��5R���[����}X��U�G�%��k~���~ݿ�c�x6�³^[�2�� �zl�롘�v������ǎ�_%e�|SӖ ��D�� ����������.=�m�#��W����d�J�x+4�r�3s�s��OVN��.�a��u7UkӅ�W|��B�0�v�zǍ��8Z��d�D��C��A��9f�u�Q��C�K �9JY��psNt���`�
G7Mc0f�gۿ㢷mM��V��S�4v͙�����M��j G^7��;�gڇ�SiV�� !K��P�Yv	ّ���l~�\|6��@��-�UPW]�ϭ��_��;`V9��I>��p⑈Vf/� 
	�G��Y���0�>�'k��ZH���EY��P�@�AA�z����xG���_��	F�1��P�Q1e���H��l[iQ'�LeݧYŉ�{������@n�<���AYҊ���8�'E��Um��J�Bop����Q_��%l���h\.�?����~�/���~�&��իZʉ�=]�������4�*�g�DH>$YY�j�R����.f��9��l��!���cD�=��a#��Ϻ�Q�-��vB�@�x�e����p���
l��8���8�\W��s�����2���M'{����_k�@4QF����I��<��7l�@or�Jł�I	n�Bkv��L���D�-k���J�w��j��v�	ZFkwy�̹�+�����5w�}ךZ}�{��oC���O~ܗ���m���G��$(�/�3����Y`�/�4��Ғ0¬1��P����p�S��~��c��W�헵�qO�51T�i�ˉ��z_G��^��`�$n��6��{������c��]h��`2�n�Ņ@����t:w��	� ~K?���
�7#��6��&_���x�=�Nt�#���3��c�~̉���_�z%�*ڱV9��_�Og�Z��X�ț�^���_
�dj��+c⮊��"|����1a�8���[!�Bѵa�d�.��5@&����Cg�K�z�Y6�#Q�e)	�%�)L@⬀����G�F��� T��#=��3��d�c��-B�"x�e�`Hf�(>�tQRZ�$��i/��o'���_�9㆗I��'rE�>���2^v�	�R�+�_��RB ���[ޟ�)�/�,��/:�E�9��i=�$�O��f��<�8��($�OX�_��pr ��Ѥ����?9r�oH��(x,&���9�
���x�K�� ��)�È�!g�ɘ~���O芀�}�qM]�=�AWQ�Ä��n���k04����=�f(I@
�|�{���!H��Ir,V���Ѱ
���KV@��d+�����(�G�7:�*�����d��d��k�@.`s��[����F`ǫy��=>���G���>z�I�8'D���^Kf����e�V��E%E�����l�bj�
P�����&0���\{o}9 گٷ;���"��UjW��\��K��o�/�®Y"�Zr��\U.��寍�+H��|':߆�ҪQ'N3Xf���m͕,���U��jJ;�h��E#jL��#��o�F��5�?n0+5;g�Z���l��Ş�n`�h^ʚô';��<"���%�A�ma�p�{�30{/-��zb��VX0(��W4�\�!l[���u�H:s��K'U��ӽ3[�T��1V�� :�������K�;D]e@x�g��ٖ��g�"�z�K��^����4�?3�)�좣$���v�rA�	��nT�1��F{�������PBH�����,���T�h�?�=L�,�ɸ*l:�IvKW?.��
�=C� �y�y��A��亽��NK���T��V*�E��0imcȗN�tMH�%��mO��=v�۬�K���DT&��5��<턞�+�.��Bw���jE���%�M��K��>��!�RNՅ�� �-�U�5nY� S�<���_��#�p_P�1&�@?�8l`��'z���+f�#)� ���dt��??���%[�%b~ �����5�˹ �̧�ɛ��g-�M�����`�6��_�Nq�KA�]%ۋ&�B�s�V�X����������э]��R��z�q7G�oM�Gۃ����0 ����	CGa�)��j�x��kAI���/L5��f��� �񾊞�T?|Oq��0w֬j���<yG��6R���cwfp_�R�
�!Y��졇�^�^�|z�{���1�d��q�X,��:-1����̀�6(��E���Ɋn/��&O\L�a^� jyX�g�dWvC��+�s|I�~@`[�Z5��g;I&�M��O=R�����G�`��'�rM��CA�Cg�t�N�E�;��4���NҦ�dh�6�U�Q�`�X>��C�/�N��}w��9v3(<,����	��=n.P8����V5m��Qn��7�$.�I%��tw
���Ĉ� q/U��P�o ��'ג���V�Hw�(���6�BQ��l#����ރ��(g6��
B�eIo#P�Ò�?�+P�Ħ���ۇ_��� ���3���p�$e�g�8��iF>�tA�(,�Q�� =� �=�����8�w���A"ДVzK���$��(�0ZT��Ikf{_υ�+;^��g�v�'�չx،�W�SLk�}<Jz�~L�rr)�5'�^朱���wi�0����ϒ� �~�MI� ��G�P��^��I�&��4QH#K�
�T��yS�W��K1&0�Pc	�R =u��(�� ҃�~��Oo*��J��%$��;?G�4�3}� X��p={�X�T���J�����1� _wB�=���8�;0��n�
�'�k{R�Q"��AFmrU��W���}���R*�G����u0�I���"����Ɩnm��.D��+��,o�y����:iR�S>�n�baX����I_ʮ,����v�$Cn]��ݏ[r1xT�x���f�I�4ߦ��;H^%�nrX� ���{y(B��~������#:�#��d6ٗ����l�I��	��K1dF�QK0C8id����E�^:�:ہ Y�Nm�(?��q|b��(�����?^i0vى�.*���g۪�+��@�=�F}z�P��4�5�_�GSJ[��w.���]Q~<N
>�+�I��Xm,ع�6p�oO�*�%�������y잴|�K��d������ER�j6�U�w�T�������1�x��{��/]���%�8�����-�T
�C�_�H:;���o�ء�B��I�{�ce��%2���g˓�-_�$��.�4�F����D�r�iG�$��ITT9^]�=�/�o:i(Ѕ����i\�Tn1�A�&���B�v�m�d��d���i�n4Lnp�8p�8o�$�έL��j2:�Y-Y-t�����U�5�!	��1153�0��L��1��x�#�i����g�c�h�9m��e�8��ǤƸ�%���9�b
����\�� R?8�%/A;�Y����$w�Kr:��w�t���cɦ������"��Ȃ���߄�rн`�o�����{��0g��J����n&�ǆ!R��IL�+���ک���Y)�]MU0��?��[�^�l[�Y�K���X�S�	�%� }�M�h}��������W�1`L/�K�59�U �������O����u}���ږ��owRU�j���Ь�gc�ecd�^R�rG>�F�SP�P�\\w�e������sH�m���Y�|�B��"Sh:��r9�!�.�S� ��V.�n�o�̋�r�nQ��k
m�o鎱(C��g�ҙ� ���G%_#��K��k�L��ż6��5 �G*�0���W�-;�#�wlv�/h����ۛ�eyr�4W�!'$��nb7�$tx�sT�ʰL߃���Tr�[���H9cGOY�wŹ#B�F�X���L�|�Iv0�$h�˽Ԋ.v�8����8\���j��Ox
��3�"Ϻo�WnѢwG��R�0����<�׮`�0n���r��y:�gxY����5�I����@!/�F�����,�yU?&)�����Qf�~.:+PЍ�}Z~��V�=S��b���`6�n��pH�5���R��KV71�4��i-јG������w^����E��689-�РLv '�)b�k- ��|��׿N���$��hG筊�Y�@7Nq3�<�^���xT��o:0�џ'�42��"6�b��_���{)�O�J"~n�
6Ƴ��qq��>L�����1���U�*�^4�:����g��m�CV=�PQ�p�ޒ#�jً`_���%f#o[��XW�y�.ss�}t(���x/���B��'= ����jڬr�D	;�t�@#����h�ډ��+��D]��
�� 0�M�#��g�������B����M]&-��z�a�j����)tA�%����,�{I�_a*A~!3b؋L���\��m;O%���'���a�vo���,��MF�����h�|
;�P�o{e:���6!-�n'�HM�f�~�P�&�`4�X�Ɔ��f��kn���@�.�n� f�pQO�/E)�`z×�����MOp��U���	�G�9�!t�&�>�v��f2M��mp .�rx����oru�{,�n�^'i�n�]�-) @67L"p_��ܻnN�	�,�1�90��	 o�z�̝6z;ń"�mv(3� ����sC�?����m��N4"�jL�.?։֔��e_I�N�<S<���^&վ�T��f�|���n��[X�V�p��f�L��W�����a��9� w��>,���.;r�W}�.zN |�R5
��?�&Q�i��T�NUr�6C�!V�\b�Q1�m'���Ө
v�eh<)c*�A�h��kh�ɣOJ
y�Akֶƥ��P-
TQ0ʗ`N�J���li����p[d�|�����E4zqf���2�u��ߐP=ا4,��mX��>9�m�R�L�n�Fo�}�*�a���z����o �Z�l�U#�� ��I��gG���J%��P��O!�gI�à�cYYKˆ�IM��т]��Ū�ɖ��i�T��"����}��G`�ܝ�wͫܫ�_��K2��=YdD�6H�V].N:�
�=��G+�bn�Bɂ��m
��yJ��/{�5l~���JK�C��-Z�6���o.ж�������Fuv	X
��-9�ܖF�S0;�xΊ�����a�oD�c��9���ȱ(��?�B�#�C와����|�4$�!��Qh@a�L�>E�֨F�\��Q�[Ann��yά��`����5q�����\�-�eD��V�����x��w`e�Y��`�Z��ذj%#Ԣ��+O�d6&Bh-y�v��3�=�eIO�r��vw�������b8ʡ����O�t�;�}),�q?�`��4�6���>0�� �q6�*S�,$���ަ���������$.(��8\��5���;�m�^�zL�d� [�D{j,\��.1�s��lR�둙���]����&b9�t�*ܱ}m�\/w����EuY~�*V�FO��4�;~���6�s���e���S���HhkE$!�)�_{�X<�.�Y�`��L�XT+b�AZ�ΐ&_�@��}���.��՝�R��XҬ��h�I���E(�(HZ}��R~�藃_d�ځ� !<����&�Y��o��r�Un���ˢ�:������� �G���!�E{}qVo�S���1'﮿�J��w��a�I����q��<�wi�!D����$FH�ҟA!8�}�0b��ş�FO���G��Y�H��|��|�?���}�gA)�q��v=<+^�_�ځ��J\�f�6�q4`�R��ϐ�R�q�#�r:�,=���ص��t�!�5�L�U�l̪�E����D�%o��z�վј($`��lQ�*}�Φ��c�A����9�Y!�ͮ�0�\S���#���AӜ89ǯ,|�����2[������?��v���?���ۺ@���_u��J�(��|xm��}�3R�77���	�����5��~����%���N ݙ� ��5\�t��O���
4����S���k��!�v��4�G�)�6���4�B�{Hҷy�D8*Q6H��ݫ`��|��Q����F�;���DH�`�:�RwD2 �r�8Цj�����q ���#Bؔ��)���5.}��F����p�x\S#{D��X�ot�S"q\�����~<�.��@�*x��2׉d�L�]����4_�Jȥ�����I�?Ța�n�@.��p~�W��\����̭ �$?=O�%$�I�	ޅ�Ez1=�w�q��X8G�Iʿ�������%�;rx�L���u��7�3-sN���	3��V�uc�EJ�=DC�蘤�WD\����6�&���������5��$���d�.QQ]J�-�rr�UN���o�*j)�1�*�e22�N�TUr�Q
����m��U
|?�j�U����	~r�k,ݎ��RTmQ�R��dy6��"��X�J�m�ʫ^I�l&�罻9_�ĵ	Fs�z�maG�巨�� !����vܶw�V��F�<�Js���"qm[�4ߋ��Nzi���0�/�нx���IG�%2�]��)��/qk�j\%�|+Gy rd\�����F�0M�4�YL��Ҷ�)Hu<ꁎ�#"��Bu=�&�qm���ak-LU��vſ��0q�Tb������8p�j>���&�ϑcW���1��D;�~ ���yF4��ĉ���M� ��o��[��)�l!��f鼞&0Y,�ΪÜu�-��c���R���.�~+,��I��r�~����b����
`ęp���KǳPV**�,�_��1<��v7�zfA)�0���|&V 3��H�|tM��ǅ�:��o~�s�Iu�͘ͅ�<~�{��Y}��C9%���ί���ɉF�|�?R��^����E�N�L��r��~�e~�5�8�+M;��M��f���1�k�Tg��辎�+|�u����Sx�8M#�%=�:�|�~6�t�ht�9N�C�m<�A	�d�#,�I���C��S&"�9Xg&��T�&YT�nh�ﺍ��R�U�~G^�3![@�e���n�̋��"_Ƭ�^�)�K�2S�*[��"����mVw)O�� TA���#���h�v�����x�\�F���)oo��X����m*f.x���o���rJ�zB �J4�.Y|OnI�c@6z����M��U�����C:H� �CMl,��~3c͑~�����j��1'7s҃^�Ir,�K�b^O!Joq3��]r��*/�p��S����u�Џ�I0�^?v{��Φ�I��E����pF�]E����Ǆ6y vS_4th��F��(b:[a�R��ˏ��b�(��󜒊ak�.2R�6�����>=��)£�
��P��'�(	*�BFC"y+�y¤���K���!P��^ɨE��n_=߆���#����@ �#B��4&�'uQ�g֞��pĎr�SRn��)��|h����*����A�:��Q|?��� 4�����{�o��(w�T;+�t8����Z��ϝI|���'8�A4u�vdu�F[K*��j�Q�̍�l+O�d Y.�2�L�ĿoL�]y��ata���Gq,���s��
��&(��
#C��G�����|�h����E-��˛'�׾�R�!�|D���<3+�0�F�+��"%�E�O]�_������"���&�1����7��^WK� �/<�Xt�F�Y.-)S�3Oi�GasV�i47��db�T��p1��� ǰGO����w�Y;�Fhi�I�C,�p�#�~�M�E,����B��y-.�X'�
���~�ݎur�(�yo��xgsQG	97yDn<?D�٥���e�mgu�8,:�T+~�9�u��_�"1@Z �گ�/�s�����A�Lߡa+�k�#f,��E�_2��jK߂S#1�|x�	��ϼ�~=��W�*�Ls&|��	�a��s������ ��})��=j1������0�-�4ּ�`dv���*�%b[FB.�*�[u�Z�멅�@����nvG����%��#��Z�p������
=��)�)�{���=;�T���]��%F�7[�?\*g��Љ�9KĐ�b�*GR�s&�֓S$��%㿯ǡ-����Ք_F���x���C�<�YWf��t��ڗ�eת8�Վ�܃���'�q�B6�Ӛ{ݖ6��Ee�a{s� gPI,C�a���[���^��W9L�����7��$ըN�ro���M��{|R�i�d�HBϷ�:7�4z�$�!�v���_U�w�	e�� ?�e.���t)�X�p4oҜk㦵�B��t�`��]�*��I�RJ'�����B���8�fZHD+��do��������5x��4��`�>��@$�����f>��n~���3�^Պ�\)ku���  {���v� �[���'�E2ٛ��t���|���H���J5�h�CS ��Q����e��������6��Q�yjm��d�"_-��'	����*�qY>��m����M��/\��u��_W��6q
d���<��FH��n����3ٯ�E�!���s������|���I����&���B���T&|��j�����9ޱ�s(���Vi#���{�֬˙�a�M����e�lS�����X@��j���.�5/�5�!e1T#b�џ!����"^5���*�� �bj��Y� 
݇R�9�}�r�Rzy�E�_�O�1$��c�z�Q�x���?��6{Y_D�K�#x:�F/]h��C��{�3���wtFX�΃xw�� ���n��7�.��i��N��Q.�_�R-���\�l?��1mm�P����_t�_�*!�X���&r���ⳳs�	�#��ܭW�����G�V�v���@w�[��U!]Se��A�����?�:��,<���.B̀�.��Z4Y�x-�o^W�����K�+{�ǉ�~��zrpVN�?��x��-�*�N,ӏF��-%�Ted�,�<���ä�̍|Tm�0dK=���P��E{ʵ-�0��K�s惿rd�W�Q���u��~��t���c�P(��K��%R
�&{5b��٨ݕ����E�ݩTc�)/gu�p���g�TF�+��]\ǅ�è$��	ˬ���>�-��׿޼;�s�!�C�ź��UފGe�@��~��t��N�a!����!�r!ݝ�8�q(~�3+K��EwD�Z�,����/]%�:�N����3,�z�n?`��O�|�Y^�Gr���Κ=c�n�Me�����s��z/��e�<{�=:�*�"��uͳ4W�~�e4�ѡ�=�&�v1a?��N��{Қ��s�a��rB�@6�$+��[��}(�����/�Ɋ��S.k-��͊���NpP���A���Y���A��H&f�A U"a��驫1�j	x�}��7V:@ĤYEt �S&<��6�iuoԦbLc��HEI`��B��um�k,��$�.���Tf�Y��f�HJ6\xrkڑY����ʖ��Eс�%/B�H%�����`�������3j�y��r���Y`�� �Zl\T�N�a� �8k�����<�a���͑�[_Y<`�0���Px'FSZX�����J#�'tv�����+��U������Ë����K)o�p����ì�>���ùk�v�fa�Qކ6\^F?�K	��N 7ov$	���+�r�6���^�B
ART�zӄ'j��]��+�b'����M~�)�%�#�xL)�h0�� }�N'����Ո���/�tE�e�]b��H�R~���V^�~p��Ϣ��X6hL��a���n���#�Mm�
=�ܻ�G���	ʴ!Κ鹮]ї�۩�#���)���}g�݋&��ez���^�;m'(h߬�.Zfi:^l����ox�?���1>pK*�F�#1-a� ��4�k�����5���uG��fɦ\�g?��q��s��E��|�|+�`Ai��*^θ������o�X{��S�{��������qR� ����A�wvTKJ��"+5��`&^]ZSa�\���_������6����7�x�Z[���r-�L$�
����y�	 ��v���8�\���v!�;~ql'(��B-0��H>��)�MFԓ>WE룸_"a�bv����J隽�B��o�����hh�I�d7x��	.�^Y!]�qD��Y��׳+K�k�n�qbO��KA���ʸ�>��]R	m����,uO�ӓl��r��4�D`.�G���m�;�OP<�z$�:T+�E�+�G꧙�~���T�ƪj����1 uX?A}z�����߿*��0K9T�F`��Ƽ/@e�_�(&�g����m�$4:����hHo��vX���A�36u�B/y�.�ϾkM]���VWD>�ڛI����F������5<��cM	dC޾(��t�
3�g%�H�⹮���d{�v��^���)X\��GӺ��ne�b�" �Wd ��B8��]�f�!��7����Wȷ\@������+�8w�V@Vy�h��G��*��g�0X�c�4�g��a5�����v�o��tӳ;�޴y�=Y���a��@pj�8��FKA�+E�,�!q�i�G^J?�J���ڐ��ǹ��h��� ����)��O��)��b����+�bM�`.�1����WF��� �a�*SGA簔�^���&D���=�	��6��V��C`�l�� �N^���eZjK�s�M�r���@��0�Ha{�Һ0%�c�߉�v/	v�yd#�"W�kq\Ov&�>ؚ��+���-��.�y��� *Vi(Ej.�xt髫�k����R����x�*9U�����U~���NQ�G����3�}��gi�ǂV�/���������j C��G�8|}��G�ۋ��!J����q���&�2 >�,�Zٝ�X(&C5��܂�*�9�mbSΆ�UG��]�="�����","(��7ܠ��������.W<�O�0݉ �#+�xZ�V��f�q��;��s�.���UD5j�)������2c�gK�Y�a\}����y���Ҧrhn������IA��R�b'ۈ�S�Xw��e��e��^��v�(_���ؼ� ���Ї���ig��V��,Ե�$�a^��#%��aU�7���8���b�/��+�(@�qU�p���S�H�*C�iW���fh�%�� � ���Cc&���:���y��-���/�N��5��%D!��B�G#�u�ݻȝ��<0�ok�y���(g�D�xN刺�kGTE�!����m��u``@�0�%D��z�4���r:5�dq��U(�&�d�A��09}�JWz�����J� �h��T@,j��"CW�@X�f۟_��������C�0��=�9��Z� �> j�W]}�{���L,b�#~.����|i��"	��G�ҟ�捁}�L���@X	�Ȕ�6�2��˞	 ��eI�O�{����k�6)��bc�6R�$>��8Y�|宁#H�n�ʗEo߱&%�O+�~.�Q��6t����ͩEKm��������r���m��9�zL�bԵ�6B��N�X�Ə�Mu��zz����(�� �H�2�+ٰ"̣Q!	�#� �\,\b��h�/�A[���?`_�p��>KfB�BٍIJ�=ScO��v��L��E���rN�,GL;}��Θͻ>W���D�q�@�	�����k�����L��@������/�����Z3)o��,�p�u-�D�HC=��wn����֏���4R�q'0Տ��FV�����������'�W��tR|��y�
Wb�@��M�K�8�2��;>t�&ʶ�2>e��T	�nz�Y�.+}��`��c餅�.���Bֳ���q�h��+Z��I7���.*�/��!7h�EH8��c�z�� �u���S���@p}a����w��̀����9���ˁ��編GNy���\� aaN��L�R�C��v�$��3��C�;;6�*�8�H����UrP�hP!�#�������6~Q��̯���~�5�,�!G���mMڣ�2�����v�%t�or٨C:M8����Q���}N	�͗��p8��a�T��>naa��xi:Fb/�졝|�>��~�H�{�$��ʀa�U]K�렂��C�,�w/qf�O����� ��}��w< �`P�����Vc鋊��~�ې���Bm� ��`&UR/�4w���[J��EA��] *��ʉ���6��byPH��ҎF��'dϜKv�^L��3eP��m�J�cgh�̩���2u�j�j���)��x�K_��\̸�كp?z��mi�H�`R0b�O3T]�v/9)��9z
������!�=��-3��SnN�����0#���@H��S}aI�ZB���BNT4ڨ]�ڵ���f�5%|��qa�l�j��2��٘:�҇'UU�}�s�O�|�r�j4&�|9GE�B�b���F��Ȧ��^}��:��^�3��������Ɣ[~#\�ֈ]�H�nW�`���8�u�T$����J�B(�RW���i<�k�f���P2a�x9���Qh#�L�brƱUy�B��Rf# ʛurhM��!�i�A!�;�V/�0��B⧁��]���2 @0�|S�������,��լfW�c�u��etD���f��g��RS
������I�[�Ț7*��S�a��i<�J�wg	�Q�K7������'f1M���Y�H<��?�)o�ߦ�p/���Z5kт�R����,���(K��Z%n��Vx�����s%���[����r�<9�Q�\�!�y=a��-��d�Vs�?(�I�տPj��g�ֶ�j���}��9�[�
f*]�����`7n�Ѳ�_�f;��6c�Rm�����c��Dz���J����A��$'�x��H��a��u�����G�{����]*�@,��U�|`�PӖ m��xPku����M;5,�<*(�Ž1E�fA)7<�A���3{ǏgD����b+?��8��-y.�U}���Ϣ�y��Z@��/R�M�_�?qh'�k�1HZ��V�zt/������I�Z
�Gp"d'��%GB^�F�i���;�=�G�&'�U��r������Ǧ��m �q�^������W�0$�b�+I��܇dM��=d	f�~�,ѓU�����U.�dɞ�CT�\��ǈ'؝�A�U��k�6���:h�����N1����`���b�w�#"1�8R]\����"+@�8D,�9z/�Ȧ	��(���U��>H�1��lS��ù\��E�I��{�L5J0b�󆭀��y�;D��o������:�r����m����*�� ڥ�|��^K(d��7-�ݬ���V#����E@P���اP���U�T{�e�S5�?��O��@��Y#|�z��PaFh�'Oɪ�8x�x��.�A�B��_>@�N�^8'�����Y/'��]ŒZ�7��Ӆ����i ��W�I��&���]6;���/�a*+D������ik<J�ֻoo��0�Q�F][iW��ԒJG�P�UN����L	�N(K寈�%�Bh��b]O_��=��*����L��`��CC��a{���c�p��P(����Ț??�����V5�Lr�W��y��mh#�	|��O����>�!	
@��'���4��4�=
�4b[��iw�Եis1�p����I|F��H7.���ٛ�="�ֱ���?�Zk[��mdq�D\�t�0���
u�)�4�
D��7k��ɟ�.Y痍�����+����.��I�5�m u�l�?}Ep���WX�M%�֫H�i�����������U�l��k��/?�� N� f��(HZ���{ �6fM���[6"`w|�-���Fޯ���	�mp��z�;:q
�hf�-̏hǿ"�����|3�e�
�`d����F�Fq>��2ܹ�&=�}��3�uZf1��;x���6�d�	�Z���S��j�Ǜ߬�����£W]h�W�<���9�����aL�4�P-�d
��õݤ�%>L[��}��[vS�O�*XX~�BG�/�Yw��˺W�j����мZP��2�:QS���^^+�]ҫ��9�(���~�g9e]#��
�里i��O=�>W�(�Ӄg@'#�W�]"jO�z��
O��A@����o��J�~r�e�]�;KW߽����{�(>���ЀJ�)F��}s4!!8��2Ҧ�J��tei�75ޱ��3(�Qr�,_Vh� ���Q�l]^��w8B'[6�%�j9��>��N;���a}ښK~�<���Rt��[Q8�#2�ֹ!�!��Ɂ��+]>�� �gA���zD2y��Ó��rM&�bX�JSB�!�B�a��=V��"+[��k\Q��a�f��W���{�-W��������WVi�sB7d]:�	�]_�Z�
�����ͮ�^�[7�E�Zy��:@ �̦��So������ݮ��h
%�뷦�}�ݍ��@���i��p��V��ay����f�X��*o�.��ldv��K���vƠ��xT�2 �6u}�!��Q�g�/�U�^�L��<3k�r %�ܕ��j�S�'mS���pD�7�CQm���c)���k�R0� +�բ%��,YllUW�����+Z#"~(�*��0������F7���$��g��`��b�]X
y�.�t���%�����ۨ2�����W��kη�r�ӂq��tatw��xA�@���S��d�פ�Qd!p&�a�U�;s&98�=Q���'L��L+�<�B���-����\�v��3i�X<]���G�Х�����d��*lhٷ���k�|E="���n,����O�".O��?H-�������;6iu�����G~�*��H��ǽ�d��V"@�DrW8$?,�shW���*�����!igµ��`�.�-�1����]b·�s�4��QZ���̾[��H��lCU��GF����&	x/�:c�d�T�w�M�����_R��_���a����I�d�Yl(��!0'��z�2�s�?�(F��ک�]H��80�l�籧Q\"�˂2�t*���;�Mk��񺅣zd�<Q��s��xDn�\�ٚޭ�s��=O�R�L)���Ò�Xhs4���0�$���Ha��I�	(�jJ�ߐ�6/���a��]�����hC���K3R�z�}^7P�Nt���]$�B	z��^m�|U'�D2&@l4��¦�XŶ��Ř��)d�T`�07Һ\l�D/�����b<h�X?�2�v�TfO����P��[jH���k�� ��j/
Zg@p<�I�x��d��V��R9�GZ�C=� �w�}[�	��dq���� =e���s��jo?8��ĭ��V�%��JfT�E�x����hH0	kk(�3��}������f8����j�i� /�Η����3n2���>2�O�xy����Q��b�>5"'y���NN����=�c�%WAi5��mHW΃ܜ��Ɓ���������4��Z��i��M���נԂ�?��;kD�TH<(-3��$���Ō��>*P�;�������d=�=�`&��Y�W2]�mC̘u�����w��!�R-C/l�������7�'�62�mcRm�ʱ�O���<��҆���DL?C��ō&ݵ����{?N��9�)��l��Y�H���輸19���kɓu�|'zn�g��I3�?Y��T��g��P��cN~���s!:ԃ��Z0[�by\�r��P	��~�j�Rx�<"o����_�2�<q%%��{kz��%>F֌;f�ۼ&UZ�M�!)��pZ^'�.��O"���bj�mhf�Sm�=a�Kw�)�4���C�A�󻭤�I3�@�N�3)�O%h�؁zX�-���X��閐KF6�' T�˵�aWzIR�ӯ�E�;ʣ>��+2�ln�H��?�-{�L��"O��:���� &n�xiuv�ia�[��a��� g� Vs'�ډ�N�x��-iTO�?U\����t<�-a{�j�����"I*�2�A�X1�OV�*{+L=����E� ����5�?�]�ͶqO,DԮ՚����� ����@q�Z���ړ��d�@�Xm3ҁA�у��_?ؒ�����Yla!���l��G�=b�j$���H��Km�A3�)M��ΆqB�s��{S�*ao��X��G*��\|1��{^�;/�F����ݥ��y6M��:��[�e|��Wo�.���~'��ͧ�I�$L>�-y�_�]k���>�1P*���A���q�*y���GU貕=�_���că'�&�?j��X������P#3�v�e�����3�?x�D��,}�z��|����J�w�s\�� 	$����7�x�J9��B�CYxeA�Ȭ��]�C�4h�)
�1- ��1XO+z�a����lk�u�fXx�Sa>��|#PšUYv_D>�oD�s�A�*脪��1���Ha��;�=1: ��#�9 ݚ��^,v-����KO��/����F�����������9���T����zן�#����oV5�y�>���q�c���	~�Ns@mΩ⓲��*�]I���g��yO�����5�j�-&Nޤ�b"V�Bd�K�3���ZZ(;~��@TK!HH�-4�I���4�N�T��_�B�������y�M���Fwn�6���|�@�M��]��y.��]`��v]��n�oL�t�[�,�.J���1]�l��R3d'ְ=d�B���i��݇�����O"�'F��L�=�`�i�PL7Y�j@����0j�10x����5)��ǜ,o|�O+�Ov=�+��M��O�.ۨJ��3��ײ��������Z��.@ξs}���F��L�؋�UOj�3�E��g��X������U��о���Ņʌ7kyUpf-70f�eHT�7�]4�7�����*A�U�p�((v|A�.�<$Jy�v��BB������cEr]��6Jw����� 
Ǜ��GD��2ɭ���Z��r���L�<�*:u�kش���rĆ�)�:@���Q����=2%M�+�s���v7����U���,�*^ /�K=F�gɊ�k�1��~۸�A
RE�����{>���bE�w#hty2��d�e���[�M�z���x	Sip�r��w���O��<�h�2���&B ��h	Z�����7"v�K���xw�>�緾�g��g*����w��Vc�6�&?D�'�@�!d��e���5�KW�|��]��]�D����WYR�,f�g��?��}B����X�
��N��9]�����SXE���V��3�����$k9��{/䉿�ÅӨƚ`�R�A﫰)X�:�al�U�TټX�j�VL9��B\?C&'ލ��'��
�<M��z��1E��/A��T�^E��k`���R�C}�ǆ(���a���|�Pj��n�}�=��L���D�����%�Ρ&i��ϸ_�?�������b?� 5(�6&�[�~	t�q�cȽ1�a31���у��* �w�yr��݅>���O"�I�S��+�A�b�?;wk�R�q��(���X��]Ǿz�GY6���W���fvh�f����D*��C��$�b�VN5_t �+�������Сش���(ԴX��%ҝ����c�)��fN��R57Y\�[En�?"56r'n��t_�F\����� �ef���rm"��v��ˬ-�/��ʊg��{3�ŗ������A�{!e�������;���;�;�a�d���T���02�N�|
�}�)
Q�W��̼��a=u$|N�,YA��sF&��\i�l<y9���5H�?Enˁ���m"s��˙�TX�8v�rhqMS���� �M�{���j�r��4����-�8G��;N7/P��z�i?�s�}}����@W/��%���R�a��Ѥ�}��z��q�fD ��QNI!��h����91�fr�z4�E���@�i��I�.F'2��sC��t��Q �-}����Vr�>7���i�t|7B	��#�!�F�Ėx����9�f�>�ǹgH����̀��������&B��m������9U�������&�{���Oۍ8B�|��>�j��U[�T�/���-��1[�i���|���)>�_�=��H��!t���Yח� E�yk=ڌ�����/SR	*[��`�֟_|�ԯ�y������4��5v�����c�+ZA�ڎ�Q�B��I�0�K�R_���SP8&�ɟ��jp�h��6�Xd������4�혃��i���E�6#�7�˧�z�� �n�sסT[��Dg�7d7��:��R�[��)���׺8L܃)����-�Vʶ��B��NI�U6�NI'p�8Ҙ��ĢON�k��>�d�K�"^CN�Vd ��������FOV�b�S��td �+/_��cNB��tENKv�+��dE����z��Y�Ik��V&�g�,���+��L��[Z/�>[
L1QA��
$�uI�j`�����d�}�)hҡo,X�����Bz�����Gۓp���0�񴑪�IL7i����9��g^L�W�;�P�ٽ%���&�����Ǧ��u�JW�hs�X\��<����u��ސ�6���Gy�XR�94����bZ�[�s1Pp:��gpc\���=ˆ)W(�Z���k�'�KA|�S*�q�oH\0@��JӤ��<�;N��p8A���%�%�����-ՒbT�/(��d�G�$C4KE���y��������g㑙f
d���~��?�*�R���%K��y�r�J�̶��7۝T��x0a��S��#��I�"*ȝ�~ݦG�+)�.���0��M��n�"�E�x=�{0:�s�1�ؘ�фY0�!�B=�O�Np��۠�$w�ͼ\x�Ӻ+��:�3�`	jb�sr�P�I,��vn�.�&����O(D�v���n�4�Ah�x�W�ϙB�K�3Qj��\xq�L���0s���՝u�隂A�*wq�$ꐃ�;�>]��9��$�_��U��v�._��e5b���Բ�R��S/￢v&��Ӿ��U�bW��E�Muv�P]���g������<b12c����F�=(iz�������^�I�Yp�ڻ�Sq��9����e�����b �+py�lZ���
܆��-b��!8��7k�&�z0��~�Al�9a�*��Z���l�U9�����#�F����W{�$�H=�BT�"�2���	�	�|u@?[?jL/���I������^����~r��!>�A`�o�j�C��3�cӸ�. ��	f8��EAWF��_�q�L��-C�'�#O!Z����Z�-��K]F(���V�e�x�!A��bﱼ���ީ�Q��;�3)	va]_������9��9�S�i��ۿXKI켘m��
�_��)f'd�baG����"�M ���pے�ʃ�<| 1��\MG�ƒ!@����6�= ��-0]6����5>ٖ���
t�{�_Bs�a1�K��y�<1m��7��Q��-ѹ+(\���n�Έte	I�YpԖ�i:һ�iL?�:�mK1�n��<r`�Ő�`��l� ��{7�mj�N�����ɍÂy��#Z���*� ɸB����K��
���Z�Ȱ�e�:�=�Sq��s{��A�		��/?@�A@��*�,���/I@������4�R,	zU}"a~���8���z���jZx,����%��U�ZD 6�f�\*C�����Hz�f_�"��y�N��@�[��,�Y�7h_�eiE	���p�^6���(J��៞��r�0�d�1�.�准��$�q�IأX����Yu���k�2�pn�J��!�$`��Vf]�����	$�f����#�DkK`;�,8��&�E<F+胗D�&{݀[�;�ˊtC#�Ig~��_�ڽ�2ђ�-)��+��΅ �_�i׮����'��=����e�3�JG1)[|M�e�i&kڠ����\dd��ײ-H�Q�ҲQn�(6c�� �[����� �n�7*y��2A�5	`jl1�pC%�-�h�@�1Zd�]j�s�=Xj��im��eEַ�R�/��oU-p�Tms��c�m <�\R9���pf�b� �7�"F|���y���3�u�s���j�i:��)�:&C�����	q��8�T��O6�\V����	/T�����䩯�u|���z����~Ŋ��8X���!%���?|�}@�ndv�Dk���Jr� *�F��`�'\�1Z+q��$��	z-�j{���_%����������TI@�ډ��Y�`�i+w�px�PvKA�g>2��� ��8C7vv��������}�������E�]��L� �H
������yѝ�hK-�T=��s]6���V�k���rH� �-S�K���S�'�(�P>Uv�[5��PQ�����r�|����I�z����ij�v�q� ڈ(2 ��t�X
R$���`6��{v[ו�;�?Q>1k�;[گqgvSX����ꛫ�yktR��o/��p� -��VGR�
r�L _ML 0�D������f�$�	�m� ��cH�����L�П��o���8s�ͺf�v��!�A�j�����hHЦ�^�Q�JCA����
|�Jٹ�I����!u�@n���2�c?eZ�l"�t���T׽a�l�@gfz����?�dh�*�f�|xB�B	��~Z$�t���z�m ��&�bÇe	��G�H��}>e�@�Dc�^r���gnZI��ȦdY�Pο��,���^��I��.G6o+�4n��&�F�#O����Ev`�
�4l�Rw$��{\b���K���7��')$��,(�J?@����^p��2ul6鑺�;�fɵ���m������j6kB���+�lZރ���6R�魲�Gf����)B�7]����?�F�q:n�ȃ�*��x���G�p�(� f]z�$x��������9���P���$j���)R�̅l���Qh�w�M'Xz�ԧ.<Α���:�����23x�%��.���6IX������������}_	$zW���5�Ł-�2�7��C��<F��t&t&L�nUK��#."3�%��y�M)4���1�"3��L�m{�j)]�q p��YB{˞�H#@h98�����&�9r��8�&�F�xbX��˽���~]��k^��y�	G�2�y���s�;�u�l�^슩o�9D<r����[�L�b�Q;;�Fz�N��~�Pbc�M׃Z�oV[G�,�t�����([$ ���@����9ɉ����yN�VƵ�"��4�2�3���"�0�aֺ�"�CW��"K�_?="Z#�}�%E������ a��ˆ~���:��EDs����	\G�;�p.
}	 =�خ���3�
u���;�n�t��|�����.���@J~��})mə��Q�C�*=-���l�J:�pMD���"�;-���<L�#��!�U�T�b
s��j��*;��T�H�x)�������}����~�	T���K���.-�B��-��I_�c��,g������:���>�!��-�L���S	>b.1�3Fn(�� ��C��I���wa[4���S~�D����
�f��-}�u�
��uI�7\jf�V�h-y���UU��~k�ٚ���B�쐩ӈ`�Y|$®�����ͤL)#ќC�逢@������>J[�^��AT	��%3��PD9���;�ikr�J�u������gPî9�-���jí~����iͺ�s��\^��H��tV������*�v$K��JaT"Y�
Z�͚��� �E£�ѫH^�=˲x�R����)"��}| p��!��a꓉�7�Q�뢬��{GHysq��۽���i+６Yi��ډ�9�ix�����XEA㊁�i9�:"�N�0�ô�k�������;�A�?�[�-!8r/�O��ҟy&n6�q�~�i��9�w����Q/ �̤��b��o�9�4�Ai�3Ň���Es���Y�h9�w��W�(��,�Y�y���.G�ަ{H��k��#�I6�K�xc3�='�_.�ZF#�ye��Ϭ�S�+�NcS���Z:Cʴq�7*���֑����A�h�Zς�l�9�=��W"8V~��ʝ7���wY����m͝^�@J>#�a<Y6q�9b��h4W/(M��e�����eP���7DU���NeT%����W!U�bR1l2s�)�Q�Kۮ��8^!߁����U��iI��o�o�ޟ�p�P#��:[Z#M�����+6;�
v���������fPQ���L
3;�"j
B�*���1�'��~^FzD��lY��9�K�3�M��0T�D�R���#"Q퀑&E+�� �<��>���h.���2O����:��ώ:��I�`�h���9
m��*�I��bu�w\�"bB��%.R��":�]e�Q�n�ͳ�\-�p��6P�á۝�JR+���gL��Z��F#�JS �hQR�Rx'J��^u�/�A1�Z�4�O�o �;Ѿ���h1<ɛg�^����9J�\��Jd����O@�O����9W�r3�;.e�6!�07E�[� )k���1n�8BW2�V�7��p,G֛�ߗh�G��ɟ���v�!t@)W[{�9�q:�z�����9v��?����E:��J����U��.;��軯Ua�)sBxX�6���Y�s���Ș�K6��mw�ݎ6ʂ
q+���-<*�#s�`|k������u�$���߽����X��<,�[e�T��:3��\/y������9�(��}1R�`����6F��ol��HH��N����:�fg�O꼘��H�ˢޱUX?�G+m�?��P..|��,��<��8��!Ɨ�C�}�jbNb������4[n3�`�x�p�E��=/�?]�8����ҝ�G�.����O��v8x�?Q�h��>�H�T�5�]n���+Fר�ͦ 9�|]M	l���������s|ҵZ�)�����g����a�9`	��.�wZƒ��Q+4|]��w~��2A@,�� Ҵ"���˦���\��av8hS�j�_���!K_���a�N��<�o�*bn*��������^��O廞� ;�w@5�b�Bs���C�{9BZB�#L��<��L�zV��\����[��e#M��'w��J
�vJ~�A&�[I���\�D�����Or\._o�R�⺭#r9�Ĳ�8Td4�{n�?n�f��js���y<�J�1���OR�sP���!H�虐���Ǭ@u�u��P�V�����mJ<���9�&���V �7�ۇ1'_KA����L/�_�_�CyD�+���h���MR�D�i��J�y)����V�hw!j�aOe!Я6dX�����gv���G��3���P�����X�3�R���ly�]�bu�'�k�6�X�Ǭ����B�W�#g�H��tU��X�+}I:3=� ��P�P����"Fȶ?c�W�*��3˦� ����j�ݣ�8�A[��m�
la=z/�o��]7�j����n$7MC��g�j3C����<mn��GKÜR�	�j"m�����j���x�A#8@@�:�_Y�-fr�l_+Īk�0m�vg�͸>Y5M@�i>u�(פ�aK=������e	I��OqL	���X��ѥ�xe,����+�������}��h��K�u:A{��@��6Nl��c��-D/Ԟ�(e�8s8��.�:������Iu�h�^ho����5�E��;x���qE^�,��ȥ�+FUN@��6�|x'�'E �J8<,H�w�}W���7��|�s�e��	Ӡ�wz5�&q���� 6���Y�tl��4�Φ�Y�
�5��Or��^oj6���|�h��vќ|���C��inQ�A��[�fї���x׶��z݆:+~M,P��|�Y-�a��;d�0�Oh��g�~o���v����j��*MNu*����D �ò�r"��bPF�}��G�;Z^�qy�w�����c5��o����ug``p��4��>>��H @�/}��1�'� Ѕ�������/����$y9�e�h��������)9��L��/� ���������?PX^U��-�dڦIܵ�s��Uhf7-K��%^}��Б�-�> #�R�e�3)��o��K�`Fhlɜ,���(0h��ul��B��{��p�-�x 6�ҦS�u'�]6I�[����SrP�����R73rw��of��NW�Y�>sJo'��j�m�C��)".��8���W!�Ɔ�zM����L?�7���S�y�9_q��	N~	TL��%�=���Z��:�ppگ�����핬!���$i$��y��ۣ?3<X��B��c�<{�� ߲�X���������1,��M�.�.J]e��g�ygc��ɣ���fU`1�� �F�w��߸�1\9��%ހ����q�-�	��D���U��K�̒O��'r���B���h7��yk�o����7��:1��2g�]�����a�Oiv��~���B!��+T?�c	9*!��`i6������_)u|���A'�!7W��:-p��^�VSi����������|�hB�V�q�:V�쟭��U��,#�  h���7�4?mu�r��3�:���(zM�{�m�ޖ3�,�*�M�Stօ/�p�
���&��{�
C����_�=�v%I��ި�@���3�G�TC:x{(���yo=�m��ǄЌtD��~/����ĺ8X��4-��������Yr�d�_��|&��x���B�[1d �'�s"�J�A,���h����(�B�k���vC�
���x���R�#�`4��3�kO
/e-qTp��R�A��uW-�����Mf��.�(F�5�����?P證�~F��`�Q$ڄ/���5,vJ�h�n�����8M�5��߲����4>z�+�I�=�g��Vy�[w���?�(�����N�N��L���\��/eGy��s��AmR�L��M�����W����	�!*r�Ui�2�e����&�����۳@�����z߷h{�OTέ����#���p��1@R��H���/�]~�{"!3hQ��8��a�Zc�3�z���'L5��=�f�����4�;�[�n�w����
����P`�_��O�o�5p��hD˔����J��������F��O?q"7.�I�/��݁4�`
��d�͢�����'��IڨvQc�)-� o�]r6��J��,�J�t�ј� �(,�%�@�t��X�▀N���J�8�>W�x��.�+��r��U�d��M �#�;�d������1�� �bW�L���n�y;H��K���i��yF�ȏ۽y�?I*�'�Ln���$���q�v�𲌁��h�!�?'m|��/E��W��}�
�5��L�2cP� ���EŇ�b��&(�9v�a!���IU���c�W|(����ͨ���[�8��B������Δ�'V!R ����L}���G
�y�I�� Yڃ��A$G���嘇9��Q�1��BFо��%���,�j����{��k���p� ~�s��2�5G���W�ЫZ�S""Q��~a� Թ ����Q8���Ui���%di�&hDP{�ɞ�Ls�l�dO�`�?}�M\�J��P1���~��2}$x�������-�=�#�Q9���K�4B���p�,Y�<�Ah ��`��y��"��\|��f��B�PBU�/JRh�o(O�:��8@�s	���{�:/B�wb_���1��A"Wg���Ò�9���yHT���+�M�7|Hj9�l� ������R�쌓���S���n�f9�J�;�j�Q��;iR[Q�.������OJ��Wr{E�C�rmV\���±[Yޞ��I�oV����B�9u��Z2R�夙�V��`	F
a4����wn�@!BD!��Գܼq��:���#[���bK���������Rg�kG�?��	e�g��>��=�A'YN=��%��mQ5��t���UF�����S������C #_�sSї�K����N��_	��C�#��m�׭z�_E3y��mݨ�|����1�C � ���k�mb5��6#��`�ڕ�����3���jݱ��vQ���9��n�Us�Z}"�Ԃ�uث�l�L��L������\�<��t��=M�`�Q��!;�
���|��"�NQ)��jY���n��1��m+#
[�"z^i�V/���s�MVO��Vu��Դ�d�8Y��g��@Y��k�8��;��7o!p�]ّ � F� o/��
Z�Y�-N?4��ŹM���(+<A
�m6�$�Mmn�cQ2�&�yX�	F�'��!��>6t�LIz��"�yf���R\g��b�˕�o���\�r���T��݇�������9�Ԏ?��_���%R���� ��x΄d~`z��#�-BH$�(l���4F��չu�mZ�K��'���$;L�W��징��oܳ�a"��)�r{`�e��h�U���4S?�V7�"�-�QO�ιg�R�s56�lJ#J}�@����@>S��0��;�Q�hz�D��-ھ�z�\�r�E����\N��B/3�7�)��-!�Hh�b!L~�	�t�@/Y' b�����8?��+�.ݽ��$�^�}A��ў����F	l�K��G,牟��g��ht���\^��ֹ#��?��x��%cT^Ze�� �|�;���ފ�E�ơNP��J-�����{��/��f@��O���B�$\�I�Y�� v&��O�������DN�-��R�B���U��3X��Ķ�"<*�� Rӯ�G��¥������Bn��P?���ߐ�P��P!��|��(���o��^�i�$�}��0�^tI�NR�����������e��$3*�I,q����	`��WS�W������v����K�q����:�k�:�L�s��/�?#�_��������1F���@ZOb>�����i'd����'�J���pXo���FS}s11)�0���O�zf��އ�@���,[�Rr}d��<�%�	ק�����I���?
D3Q���֡H���-ra�e���-FveT�BI�9�E�����b�0��.�~�ty�����B��C�[�[��p�)0����u�S��o�@��5A�ĝ���,�,�xs�,zą�i}@_���N��m �邡�x�9��{���C�rȼ�PߏI\�`���zsv2TM!Rz�_K	D>+ȧ���uF*�*L?*V��Z�b�@_�h��zh�U��-�➅�tsojW�B����k� ��$�}�ƦYN��[��O=8�!r����$h�2�a+���O�n�����\-R��,J�\���w�ӀO��A���.Yq�OZO�EGZ�ʢ�f�Ǜ������+�=�{�&��N��B1��j���\\��;���Gj ��݂oi�8˞3�0	����*}"�<�G5�2��� ($�˻@uvMܜ��]/�_���J�� ��GMN=��Rj��L�l0ZxGo�T����gnI(�z`S���Q�xR�@���x^��F��� �|��; �����]a�-H�ט��!��-�E��ز����ȁ9F���QD6!D�A��3\�����Ѐ��-UI�bk��@4�qK�k�!�YC�-�!���ꊃ��xL�नqF��m\HgѰ����	!��P�+1)�����<\'�)��XF8��2B�d��n�`��Q�ȟ���7CJ@Ok{Бe4;�����HƨJ"؅?��Q�3��J��_���\�������7U>@F�64��2�(�>�3���mqķ.Xtp�iً8�$�#-ī�.$5P �t��=T��h����%��.�#U��T��oL�������vL�*��jG�!�й%B���u ���@�֎�(9�ر�����.X�L\���5^S��/��H���J���5M����HA��W��Y,ω>���C��
G�Mn�|ڛ�a�kT�(ǽ�1�d�mx�S �1�ZP  ��x͜��;�K
H��K��x�si�~*��@hU�R\7:0����͂gG���ф�`K�M�s��hw�F탣bB�h|���L��Q�ҏ�r�u�<P���C�
{,�4�2���v��Ϫ�|�^��ti��=���
J2ܙY��Ə�:{[5ɍh���Z�����2Y�A��K���9�[0�=�w�<���A�c��5H���Ն��Zuo�O��*=��O�I����JT�X��'qJk;���3{�i�n�	��F����4Mu����ðKJK�;�>��쾝����m��S@�efH��~�&~�����iQ�V��k~�9z�w�l������@7�F��L2����x�.�>a��2�t��xҬ�>�A==��WlB3B��_ ����꾭c"jH~� �� @����:k������*9��+=�3ѼU�8U�3U`�!RY̿͢����b��	w�|^��E���0�-��ຓ�1L~^����?b�x����!/���=��;,�r]��Чe��Tu���?Ƞְ*[��!�P"�Wv��-�}a��(U�犨ײq0�=$��}L�c.S��׼
��O3R������:��܃��G�d�|QMט�c�U1n1NH�+2"���o7I��k����}g���k3���:ga!�`��̱@�۪�]��d��F�^��%��\1�_��1�w�%5�a_���z��5re����:��	�g+sO��pjР-ȶ�<pZ�ww���g����b$λ~���y yMo%(��lF���"�Z`�$��V������@��;���L y��1(+�l�X1,8�w*)�H�Su��4@g��W�g���8��2��W:���$�<�I�q�QZ��n���	�Ӌҽ֮Ԣ�� U����4��4�`|CC��u�14K��M�҃�8�T@�\˵b$Y���q��A��\�nUˌz�=p.XĻ��ث�x�`��Ovr�_��fN/N�F�qn_�M't|f�v�6W~����SUFͫ���5�X��a@��4C[�Q^x`��5i�������|���K���Ze׫�"^�I,���,����q/jW���[%�L~��!=a�!m"�y��3$�7��>����x�iy��|�k�k�4�u$�e���֑qO��b(c���h�24MΧ���Sm6���dW��8[��1ϷQ��^08�,�Q}�0�7��=�(V��I��cָ�B	r�����!����|��,7 Nr��>7�m�^�S1t5#����@���[4~��|��UN��  �UXM�����QW�)+�ryo���[}�U=	�Ս���c��_#���)�	G�7���M�T��zt��q/�+�O���"Qa��lz	w)vaZ�Uv@-�zr�J���X��@�$	�����w��s�=E/��X�ҍ��sl���3��f��hYvuF^�ÉR�C\�`�LGx������4��̃1���u��^��I�� ?A��^
�8����%qd؄�o%;@����E�al��c�d�p$�!���c		�O�+ !�����k��s�޷ ؇��j�^?2�3��h[D�P��&���O �̴-�S'J+���K,^�{�$@GT�1ipZ��yy�1+t6����<$�+�!K���QTgLZ���
jz�x0~8���������j E%b��W�lϯ��z��O%�S�l t�� FD�$Qz�����(=~#�z�g	'm%�W<�8�A1)v���}-_K���*z#@�+e	z��583�k���h�1$L;q�Y��p���=e@�?�)k���zŭ��EuH�n�,_��,'9&��a�_s������h����U�K�K�x�aB�<8��3\rn�i� \2R�����uK�m�1�긫G"G���*��n�2��Y?�o[_^
�#U�lڷ���~�@
Opܯ��Z_S��V��T(�0K�������S�GAA^I#����Fjy���j9I�D��5╧:3�@�E��S�q&�&��.E��n�dԔ�@���G��YU�cp��;���kH�yЧ�3U�N�J�?mJ9�V'`i��ɪ:,z��n��z�DXrO����������6&L����,zޛTj����>�x�v�!���m��=���ΰ�T(^�B3�JO�z>d���'̣]�l��h��y�l5�3�:&�0��h;[wmh��c��zI�Ve�J�x��)�5�D��ټR�$�EZsT��UP6d�W��I�\��B$��`� ��ճg��-�^v�l��!�(�B6P]/TG�TڱvN;�f��|x��Y�ݹ�=Ɨ�i���y��]C����=2����93�U�
������� ��D1��#�ގ��&����R�4GIV�D� !	������n���LW��k<���k�>�mn�)��d���tuOR��߯75�1?iD��d� �` l��<�e�ׅw<*�cjy�wǒ��QJ�4A��ެ�]WV�2'K�Q\ki`IjUd�X�#u�W���l�颫�17D�۝���Q��6�&���>����+��h�[+R�}\�8L-@0
#�n���g��V?~���x�1Ut�@����/2�
y���O�f���=WVs??��K��b��WE�9	ۆ��1�.���,���YJ���Nmփ�:g��fY��B�M�����ހJ�h�7�^��2�O��'&q�or�Љ���A��;��!�]��f�冧�X^��Xp��������y�&�6�����]X�/�O�y`���m�J�E�����w-���.�F�z�5�+��v꿌Q�;,M=�\>11�dQ���JH$���
��n%�^�|����+"Mzd�u=�K�Ȗ-�Nj`{	{���N|iE���Q��K�V0�:]�t�
|�����P'��\Jn���qv�_��e�M����KV�._6�l��?k_�0z�t��51=��59Gˍ�|�@�5B߯p�{y[��j���xٯJ� K�
�h�Q����oq9��шX���:�"�9V��eo ��9%/vX{���pO�@�B}bU���ebqO�xc[��|����lٮ�`���u��h��6�ҡY�v
Tàl�Z�������z��g�Ϸa��w��U�È6Gɛ���(x�m�_I�Nw�����T}���`]�UP�̤�$,��JX�p���o�Ņ=f*��m~߸Za���%�����r'��E�V���j��˼�8�e,<*��� :��W@S�3������&\�g�q|{� ۀj���\l(g�6��p.8�6G݊{ĤnZYf�Ly�4o4�H F��e?�b��O�		�@v�<�i��r=w���S�o���3B�Xhj`�ܖ��}�ۥW�ے%A)k �W��X�Ȭ{�; e���Z8��cs���Q�� ��=X���Y^���AV��,x��З�`�t��0F(���)6}p����S:殢���1E�e�8ǯ0���Z��[��M����ʕ`��E�%����e��Z��Y*�VCI=�������6� ���c��H��+���p��>��K����&cޜ#h�-��g�F���N���Tp?Xo?~ 5��:��;;!�Ar��'��id@�G'����ҙ�^ij�X�n�ӧ<��Gr't2B�@5��y��S�,�N\[�p���a�c���p{/�X�*UT�S��O!�C�$���`��U#ڲ�r��(��a��-�+�!��Wq�����Ƿ�����
��������A��`�U}���Hi��3���φ�=ǹ ?jq�/D��$�t�-��|6��䡌�Ε~�U� 6�A�H"�����{��t%l��_4f�H��{ЀI�n��=1^�ӝ�8(�
J��ɗl����c-}�=�g�>�/(�(��E�Ԣ^&iiL�v�l�I/���9���p6��k�����,NO<�c��Բܿ�aO�>������o�c�p�[-ڀ{�J9��h���gq�=�뒼|a���ļ��Du��_����I�S5u��0�C�C���[g��{̦�=~�r��ȦP�jM�����P	��q��X��q��=@Y�/ ����[�V%��*����������1�Y���86��K�F2��9B�Y��ʐ2��>��|o��'(����R��30���/˽��'�jZ�ŨnaVY]�We	<9�7@=5�6�PWp�k-sԾ`L�)��CРD�lZǹ�[��6mz�鵺�J�ŶJη���?��G�s8�h;#��臉��	�'+Nci݇�aG���H��p�Ҋ����͟z�������a�����
��b���
e���@m�=�9F��4PϢ��������\�v�\I�407{eH䕧��:�ԇ���x��k��7t����3N?M �M��"���`X�ᦠ�(V���y�n@�t�^��xL�UZ��;�|�O����ݜ���k����*;�dέu�N��ף�ZR�1�gFТkf(�G'n
�7��ȷֹ��2b6ll��jS�""�J���&��c���YhW���p;җ��Q(z�1_3г:���$�Q|k�n�j�ŒI�����+)�f�Kf�`?&W0A��R��TL�yyd�F�x<���t���c��w�$�r��<=��9)'~�C}���!���`Y��?�D��TO"�Ɠ"�I&�ˏ
��f��+��ds����MJU��P�ԛkP�M��5��A��d����q]��Ң���li��]�bx��[m}��Rá���&��� ��L�DlTP�_ɣ������>��s&�;fIMO���ʵ�����o�����`���5f��;-l{0>F��c;�1 ]��f�%H���ђ��</W��=�KM5���%�f֛�k´(�<r��P�,�U/�=)\4)],��g�b�
aĥ�|������iU-~��M��*i���a��_�g�S�j<�_s|�w�H���!�K�o}�r8�T,ۊ�m�p��]��=�@ef<�C, Yx���R�T��?J)%�Al�y���f���-,�H�']\x[*��[� y�m��4@�@�RD���o�k�C\��f��)���G4�������Z��[�q�4���;?�Q�l_���Fm"�<+/H��̲��ō�3ճ:seҤ�礢a��W-�/��S�Y��,�ɮ�Mӆ߮��:H��ʦ��/����/V�dG�t�w]]"<N��%��������.�ό�Ġߨm�b���C떘+�0��G���=ǎ_Ze�x2f�¹�q4/]y�3�]����M^��}���K���UB�R;��"�1SXT{���~����6,�������S6�c>��裆�j�����G��:����_�KPR�W��_�u�~�Sʊ������6�o>�e���R�/�Wϳ��0Q���ȫ/���V�`��ys��v�L���&[xg��(^��l��,� 2;��\�=��f���º8A��BvXe�gje��F�3�W}f=Q�@��p���RG���u�6ɝz�Z��I!����Eѷj��w�@C$������*Dl�v�H�'������T��,U��\P~e�B�vy�N ��F$������r�C��a�����6L��� oQN�Y��������#�����Y����k��Գ#d�4�eG����B���٬�'�<�	
>�aH��L{|w�Kk:�ݔ�`MF'��tuC�@��:��HY�`(��2J~� J�Qd�:�����^h�=G8>J��}k3 �?�*N� Ѓ��P_A��i�A{?�F���d�;��y�С�9�Hi|N�A�����[�Q$ 6�W����'����^K�vi��Q���+��}�>Q��� ж��@Wi( ;7��8���J���3��+ײ�G�]���m�Wt����
낶�A��T8y�)�]7�0��?�@J���$i�9���=�*MIܸ5���-ls�^���G�lUm��@O�B�~V%ڨO�l�.&�Z.*�
%BT$
��K���n�c���H7��D��A�z�̝��{=�АU�x��QJ�Z��q#�ڌ��}�-ɸ���CϜ���� ��~�[sD�7ˌ./��zJ:F'�:d�M�u��LV��^	Ę%n"7��5ef���BF?Eߛ*���9��,�G�f�I�D~���ӥ�3�u��i��Iֳ�.�[�2�0�t�W9��65��jU�.���]����$EUu�&55��z���0�d*,:��}��>�x7�T��V�����k0I�	C�G��e�	���+��go-�<� ���-��¥�@c�[�F��z$(@�F��]�6��k@,�<���(�欁mIo8&�"%L*��t�4�|$��+��u��^.0���T8�8�*��gR6�>��|�+��:5B��F/	�.h�p������U׺�K�oT�~d������~<�3z���۴jK�����4�����'��E]v��������2�G������Ĕb&�/�Y+�0�E�=-Ҝ���]�����Ǡk����t=?�2�[�L��mZ,��9� &�9�.f²��ϬX\��Ep��nd\=i�v��¤5pZĮw$!��5�UO:7w���t�
��eT��ng��&�Hd������C�,0g��ꂴ����}s���␪wn�+�cÔ�k�_���6�'=\%���o߀�#9:�ͦ����<��;�P<��F��iB�dht���O���szM䯼xn�b��&PM����ՙ���?[�ٲ��(r�F�)���	,0䅒��O`[�K����4�~�#;�L�������-�S3��d���������$L`�Q������ڗT����J~&xgK����{�&��|WI%U��3_oC?�ֻ�%W2���az����ŷ�Be�o#�_{�HXW��	a��dA PQ�5�*A�^.'%�^������l�"�-��QQV�68˗F��r��m��m�Ϻ/
0�ax	"�bD��o��z6�����>g���GE~�[��B����T؃ǹo��S!�ݐ]}�٢lɽ�/ԝ.��XudzE5QY˭vTa�IǪ~	:��"���/u��gi:&�(c�s�y��5@%	�p9�9�z�(T���xA�zq��q��e��1*�J�^Pu3����j��d���� ��w �/"o�_;�¦kO7OXP�/?޷y��~�ԴR�=$�gd.�2-�Qr}�oY�?y��i�>3T�WL�O�g!Кǭg�=+ߔ;q�D�?ܮ��@!0R*|r����������Z���`TE�E�G��{m?1����TW��'����@��i��sLț^��Ϯ���@�/�R��H̴旄:x�M@u��F������zy.�"�J�@]�����
G$��?M�vV� ����1v$2nk*��X[��Be�?i�����>>۹W�)1� ��LY��Ɛ�o�0-�����U��ƕ�����}����N�MG����$����w�%��/��re�����vV�G8�|�c�-��]��?�IY��
���'wP�p
���� ��jD7\���O�y�J�"�@�� ȵgD�K��|ܛ�4���TT7�a-�J"[�+
!Q�y�z�
9�L9�@D����[�'	�lws�{+��2� ���J ܐ���Y;I�!�"��$UB�VE�)�A̫�V��Lǒ��e��>�*���Cn��<q�V�7�TBX�!�񺃘j��ʿfWM#����*��R��T@X�>.�����w��K&cC�~���aB�3]l����ܴ:�݀�N����M�!%U{�5�	��-_C&��D�R5���1#�K3�b|�6��L'+M�EЁȎ��S�@���3x�T?�w��,�&�n����c�S�G���=͊0��;"o���	��T8���
%�!�n�Q����h��J2������õ��;�]� ��OLwY4Р��B����_�����P���F���n��X�̻�o�I������D�a��	�Aaϰ�Ջ79���jZ"~�\�V�FNQ�y�a�q���F1�9Z�8Än�ؐX��� p�$;����ULeFk� ���X�Lz
3p-ҽ�\��¶�1Pr��Z�eC��z��G��c�	�\q!2i!'��n}~�rex���`��,e"�a�Sস$Y�zX�ZvS��[d�s�r�;s2����i9�jwٔ���f�ɤ�'��kZKn]�2�h۩���@�"�k��Bj˙�'�^hu�ت4}����3�A��y��5{C((��Q�Ωsc���%��,�@s��"��".
V����b��~��e��\�Ӊ	���>k#[��A��ʇi��Rc����izq��}�D_�{u0aS��E�-���ق
�o���pn|l�a?�&8��a�����ٖ_�e9#���	�Z��,�=�����l�:x�jw.Ay#L�T��i�{O$���q�`��Hog�����<{�������G)6�
U���H��s�N�F�Y0 �G�&��Z��=�N���k����*]i;��Ѿ�鞲K}R'"RSWB�]���l�05���w$\��C�M���a���*c�x�]��2>��:{��}$O?T@[�Y�l��`Ǎ��/Ke4�68�8VY^�{�=F:�M���⩩~��fM'�\I{�f��h@�]҅������v<�"S���e�$>SI����/�o�>��O`�ve��M��Zu	�&�~x�{��;I��/��l�X�UB۽���}S��?��kS�,�.M4ϟ�6� ��+a�̅� ���/�c8,����]&��ۚ���4]�	a��b9�Y�)n�׏���P,�<�S�
�����&�{�M7'W�ǂ߯sQ�Y&O���c�������O��LA�6p"�U�'o� ��ٳSi��h���u� #S�oB��5O�$����I7�k���O�8�	�n���=?_�X���Xy)�GG����	���)�70,���G��ȵ��}QH��I1L�j��� &����b���ҳ�@��yܶUNF��˸�E1��=��%�?\��s�0��I�S�-�o����*� !}�ko��α��y���.?�ɖ�)q��M����QF�#4n�ۖ���/З�w@X�a-ẗ�P
#'�_|�%�ń>��\Yt����m��tǗk��oj�˲�AR��<��4ۣ~��qSy����˶ɢj�xl�",�0.���h��d�"�y���V�/{�,�x�O��������Z���ۻ������P�L�O�&���NXLh?�O<�����$l�)�n���..Ou� D�~�X�k��V�p.ێ�C��}F=��ʔ���cVW��ŝ_�h�K\۲���֦�c*�"S���6��y���N�эdh��d@9�j"�M;�N���ҚۻuW_��<����$F�tA�sm�gۖ�Uo�ٹn�jᜢ������0j��QS�H�w�������p;�%��\\�����X	�"���ƿ��K���yS̡<�S�7�o�J��QӎЖ��J9�lk ~'�@6�bZ8z�օ�+Fl0�9o����^� ��FՂ�-��lU:l�M;yf��}�E�������r�@?}V��b����z���0��y�ep��o�v�j��Tߚ��V�(�;/X�Sp$Ţ>G�Ǫ�P��Jm]+�^�8h��;����aC�x����1��n�B�#l%tE�LGH�3�iA�X�W�{�<��Ľ�O�2}k���+���ұ�;0��!��D�~��\������2���t Gg�5����a��d��I�;�L�}"�u��)R���l�(����>�`�#\���8<&~c^��r�ǋ�)߶�����}hX>�>��IS����S����Z=�y�x���3�|0��ǆ/�M�m��k�f��}�F>y;m��;_d+f��1�3~3$q���p���Da�<F�>�p��AWs^���V��d~Q#yuP��w	d?�u=��H�}�x�w�_�V����k�\�Z�V��9�����ahkGU�.�� ���F��x��5�/s�ja}�/����� �Qs�Zف�$�.���.�Ē��M�ԕ'u�vj�췴��2�j��o�K�=a}&ݐ��s��{Hf͂��:�.#����[����ɛCD��9Jϱ
�yoB�	�%��p�t֙�*E��˦1Ϡ��-�*=B�H�!Vq�/#v:d� 7�GAf�,�G�|	5}�m<~_%���P���kI:s�ԯ���^9;��7G>Ȩ�"�~0:��N���jD�st[!6!Q�a.%ki�VR#ĸ��];+��ar��g!SGZ�>Ü�mg��� ���l��D��G�#�3r��?{]�w<��c�>X��a��m�O�������R�
��9i�׍#���O۩X��7��Zy�"�|z���Q@����1Y8A�����;�����1���������{p��v�c�s�MB$�\w��]�3�\�%��G;��G`�b�Q%$6�Lhb��}������;d���y1byɼ ����Z�W
�mG�7�p$f��~�C^����S��+-��9F��l�儥�np��O���K���v�ˮ�-<�VG}	�Z�i�[���=��o�1WГ_�ǅ!���u{�ڹߘ~0�^]gQ�q��jC�(�.�|G��7!�]eQ]o�����p����L����dz�,�7�8�g�~q��U㸰G��|m��G��	�@t�8�~ת�&������[���8�ZZ⋤�dDy ��R^���t�om��9����CVn��2>��n (}�/}ў�2����Z"�G�x�s���(�S����߲;.aP2��P"x}h͇{�'A�&n��v,�_�^���;������X�Ϝ�Âz���	j�h���jq��n�(���t�c�Aq���9���eS���������,��/����qa�T�ȣǔKQ�y>B�CȮ�U(=���'�/V���X�:�߷U'�Z�~W}m���R�)['��!��02�EϰΨ������@s�s�o�3��2���g��c][�x0)���Z����_�9���by��F��V�m?��'��іG�M��	��:��H\F�1I_�<)ؿ%�~��j^!:�h2ĪV.P񨭙H$������$����p�%��w=��Ӂ<����A !AGK.��KVN95��pEƏ�r;ڲpx	凍�q:�:�G9ū�|��+��%�3A��2�B�t��(�D1��;g7ۛ1j]�	�������!zٯN������펬� ]̶Pr�O��=�[z4[�g��S�ϲ�G�}��ދ`eX���-�uF�d1-7��ن��|�r� ��u�u��I�3-8ũ���ȓ�Tx�	Xظ~���b ��]
��[}�A���i��a=���;��nlȩ�����`������>�Y�" ���Z���1<�1��BX6o�Jru��2��6d8�B���*᪦�5.�S�愷�A�0��cZ����̊���}�D���0'�q_C?/6��=@}�	�B��r����Tn�=���5_�Z�(��'�%�.F�]F*���?ɾ�M_k�~�?�F�����<I�I�אb�)C-w��6U���v��%G��S{K8��E�*����o��P�2�y�9�u�5���4!]��/�0r�_U>��C�g�jşi��=%X	l{]ܒ>4�����bL:"��2(����s"�bw�=ƺ��SUD��lQK��3��Z��V����K��ɞT1��u�uO�� ��0QsA���{8QP�T�s1
sΦ�+6�!�����>X���K������CT{
6��=n�s��o���7&&y O��H}<�����T^N�#�}>�?�U�	�m���6�=���f$�����Ѿ�������$L`c+�w����I��SC2�cbh`˰��2�l#��˄�X�*�R�o$�_�YI��o�˭82���A�E��ܥV&��=�����.Xi�++�@�WO���$�ݍ��Q��Z���.kej�E� M�b�!i��j�1�$�� �����Q��֬�P���.�}*|��X����E}���i�R�I~6`����J��I���x�*Y։pMJM v}�⢻��7n��'��>��C�ص��m`��~/�M@��39��$[yܨP�2x��5������D*<� 1P�L��ixZ��������S6�m��z�ٟ����C�+�ۘ��B�5R'�&��P��B�œwr����u�s�eI?��@?�@�㰾�g�DK�Q����!�3�v�8��Q�ovS�n!���g�_À�f��6/����$%�G8hJw���$�p!1s8�n�ɺ�vK�-���
SΕ�?9�ܙ�x�x��.��!.'�H�ͅ����`v>YH8)T��+ɹ(M�˹:�y�ɠ
���t�|��A�wJ�Q�<�( ���sk�N��C�a��pO�w]�`����ɻtF��L�x��o���+;���W{����ϝ��%(Q���<�,�����r&&z�1+PS������f�/o����(H���a�^B�	�,k�j��$E�a��<K���m%��Yt����@U�!�`��j����c�ʺ��[�okcʒi��Vh��M�|��E�|)����U%"�D6@ _mU��+�[l��z-�e�v��ý�8G�`<HK�4�J峈��8���a�i�#��$��X��K��AjS�Q!5.�� ~�xin|u��N���m=�C���b�[ձ��#��s��狜x��r����DE��3��B]�d��d\dӜsTn)�z��D��}6�i� 	���F�yS���U]��Q���-�eC��?�i�,Ե���70�I�uSm�]��݋Ef1��A���%�:���ŲB��� �`���z|�o�?��-�؀ow��i���U�2���->��Xng!ǋ���,
����ZJ$�)�[�f����!�3��#y���0�I�@�AO����Q'xN����ٯELP��yQ�[c�[����<�%��0���ɯ�8�Ak�h\����Ltj�b����\l9�a6jo�\�^���ֺc��S�6E#ʋ_X��A�Ш�L��hh�/�A�Xh*�s3t��� :ˬSr���vhL*Cn��=�k�%����8�^��S����uqs*��;�<?2�s����(n͎�[x�aw��D/��H�r� &���_='������$�`}�#�mV`
l�U��RH,#+���r��{���0�A�G;2]�t��\���-��.��8��k]�KG\-*�i�~���PD�����68�Ǆe�ƖR��2y�M��0�R�wM��*.�L�Ӿ������ƭ�F�$�����ģ�J�uzX�$�ȈAr�)0.Jz�w큗P$�M�JP�ľ��o<!X�ݒ���&�	d��Ij���ӏ���[�W����\���!��ª����	- JZp�w���\Џxܳi�������b�d��	`"8��~K�BHD�Gŧ�k�T8��w۲���'�_��Ҹ	v�(��.J.!�h6u���Eog�a�Gp� P_S5���HgS�v��1�ރk� �
g,z�M��m�`�#[�uDoЛ��u|6\6�	���@��F�>�?	1`*PE�b`�H����@����5��f����S5Q�0xZ�9]�{0����S��	H6�XZ�;<	��b���KKn:δ�� �G^��%��ltP ��}�ˎ�܋/��f�v����|��͑Nf4cP}�:�W���1�~�h�H�00˻Sl���n�Ƥx:I�t<�#yFAM\��=�u-�H��z�I����H�9���)��[*Z����C�~�[g��!���Mb`5*���Y��S��6�sw}��j沶a��!4����/��[3N ��i�s�@��v��(p#����H�,�	r�����4��)�73����<��
�5���}�&3N� �2|��dL��P�n�)��M�d�Õ��j4W=/�kа灮���*�'j�1��J�3/����_Uq�[Mb�5+��U�]A�[��!���$�~��%/t�����j�����q\S��uH!�m��V|/?ޡ�̿�P�G�����+HKw���l�Ngj[��k��V��H��̝��`��R[%��T�;�ߔ�a�<ő�s�D&�w+�7�Ac����M	҃,�$��~���͕|�L��n�~���&���Z%%(a��Y�a�{���&ݑ����I���/��a�'�D�����ѕC��]�G]��v�>h��Cs�9���20;�}��I��i����FA�'�>_� ��������6�Ujm����;׮�G �����jI���I�GU�i����>,��XMp��0�!j}~`oBy{�/ڎާ&O<��`H���F��q��la�{����ִ7�3�ID��1?! :k�H��[���0�r�g�U���)�y^����6�9�Yg=ޝM3��^޷=�q�8��.HYi�s�͉_���pE�CZ���miW������ݚ�QtDw�rS��@�>��F+2�Itu�\3������t�'u/����*h'�Bނ���е�l��>�0��(+VC����~F��l�η&�*L��t�Hb�'6ۆ��������[%�į>��u�����A2��p%s�n�ώ<s�:^$�;��3$�ʡK��|I9��Nũ���e���43f�������s�0�b�-TP�_���a�ea�D�8�����ٽ�px%0p��s2�M���n���o�<�F�՛k5�o�7l|ؾ�hp%M�/�X�~�o�i�4�)_��<�{�h��yT���-�x���4�Dc�2E�t���ڑ��R����Z|�����z���8�20��
'�����0�S�XԿ�����R����K��PB׌x���=��wG�%�=��Q��ƙo�$�<��璜�L]�a�����N	�^��Aq����WM�#��{!=~J�0�
����O�S�"�ϵ��e���EJP�t�u��^�/�d�pvsh�e��7�88���&�'2E�W�Y*.X�[���7�N��Uf���cV�1���]9b`���"����|�=u"R6$?5\�9�>�aYz�]!�CY���!x�It��S��r�����z�/{������`Dx���r%��p�:��@�ߗ:r)3tF,�%�H������>��;�YG�I���G%J�y��7lG#;����Ҍ�Ge�wP�D�k�ь�R9Z��4�[^���6|�"кF�8�p	6�l�ъ���D:C���(�]�lh�q�=��z%a�*UFq���*"�c��w���1 �k��"��p�~j�e��*}�#�������/����8��y:�����C�j����[��q��hȅMq�m`�+m�~��],T<i�	˗�� w7�.��NF�!S��P����b�+�	��4��ڦ()D�2�AuC8�؛y&��V$�7_ф�LN�i���@��-r�C�\G��'�/xt��Ι/t#]
�X)����Y������~ߴ :�\aW]'q����#�Z�\��|n����˨�Us�D���ع�q�ڽ�Z��|�wr*Pk0&f�+&!N.mm� sh�-zڢ7j=^<	���&�Uh��̒�MV��ĳ�>$��/��'�8��^��q>~�t������7h��p�tz�|���:J ��7!ͬ��ޢ�k�sV�7-�
����k��߱��|\B-�aw\-3e��˵�I�}��7�zQ#�ӑ�)��:mF�-ߔ�rжQ�̬�P#Ȩ}/�R�l7�2��r�����p=/Ƒ�Uj�z��}�:��Dvy�����ɥ족J�B�/e뢭]�`��E(Y �/�[ƙ��G5�6#L�N��*��y`�Ũlڣ,7��8L���
%o ��������.��6k�τk#ݾ��E9��i����L�i���K��M�]?����~?V�x�:]V�*���'����68NQ�x����D�-J�4�y��jkf���=��mK �h�z�N��w�v����/���mR=�6�@$��y��{��#����$� 𺌓K�$��/�v��[� �JBu'D�H2|{рx'ޜ��M�������V\
��!����0�ݐ�7�ǟU�n�w��]���T��*z�u;Xvsc���[ԃ;{�lO_�?��q�)��n�]�1��XD�[���}���|ր� P��/6款���p�� l!x��I���t�.�O���M�v����l�ݖ�DD+�(�Iu�c����[9��=��0�+��G��[�lc�$AJ�9x_8�<�֨��-�ۤ� �jl�>`^��׳��h�����E�[,�ܜxr��T�P�!����U=ui� �~Yd����	Ǭ��i#�"JZ����W:���D
���\i��>rt:f���&�'��3�D2 X�Yg�y�󽺾~��Xt9[6+��J�ru��Y\KӁ�cB���I��cd+^�a�+�}F�
�^�c�P.�����8��7��]��p8P%�II f�o�>:�H]z���B���igڈv��Uȶ[�@������K�Ǒ�g���K�_��_�։���,8�v���u$/�[##�~�+�_�j����U��w��eF�
_� �R4<�V[*�9�f�W7���l!z����qϣՙ�u��Y��5����+���\E~v+8�6� ��!w����yŕ��=�
(b�>���:7�����6h�2 g�'"nQ
F�(��G;:�X�>NL�?\J����^��T�GbX��E��r��CӿP=���[�����Y�Nr�wê�M�'��3�*�?e��YH�� z�,���\���m�9�k2�m�C*��4i0$��YFC�i"�2��Z{��i	-z�G	�laT`Ň+�|�1�1�O* ?�Җ	�m��Gxq<�9V@����v't|�B�=��w˼}ᩡ"���5�p�WޕLpY��a��7*�dh���A:� e�Gq��gw0�t�v�q�)4~f̰ƭ�B�,��;��h_`���L�j�WW2�?�Pw�]�D��U�.�v�'cɏ�ԟ(@�z7�Q��_�y2ڨ����i���»���C!Qu��h�SW
��w���B�lj�>L�
�O� ��O�4��>�myF��B��w��A�{����@��\���D�z��&���C�Z��F5����z�~��`�RL��v�W#a}:��� i�����e�Աn"�����U��6s�B�0��熐+��e����* y ���7�mhN{�ii��ckuJ���g%e���QAk�M5Xm�b�"��!2B�3%`��M�BF��x>���#��;���!���I�̌^��ksꂥ}ɘ�z�X��^z�T�`���v�j�i�)c�;fQ/�ZMƀ��򙙾/]�\��$J�mX'����ã�|�,鵶ˇ��o����O��gA��f�����y3���z�5״��>bC���,=j�y%��'��v�K�z�X�a�f�Q���I\DY�T@�W:��Ld{0)�:�r��E�#U6+��
ֿ�W{ջ�ۅ+�y�!g.�-�X��U;�z��ϸ���|ø1��B�fS�{�0`��Q���&c�
�H��V�Ng���@����g=؍?��w�����P�$�@J�D���1��g�c=���ҁ���Ee�,ǴҠ��F���is�Uזt�HY:
��������fi��e<p{GzK�Ґ����{�c�K���Gr|��Z�w�9�
y�l��>;�v}7���r)��W^�e�{x�[��_����GpJ�~+&���r����c��q8�����ʇ	�w�yC��G@��T���̝p��J�1�K3l �c)�;���	�%����i�­�Y�:��Լ�a�5%S�&���Un���u��F�B�'�b� ��Nu������1�B+�tV�����/db��C2�l��{����T6]�.�ꁥ�4T�����c�G�O�m�0���HGJ�(v}0xqqPWv�����͙��ֈO̣�������.��K��2�%���CѬ�M��ĈL��Y��E�'��r�#���2*S5~�Km�e���E�g�5}A���$��f|�9e��=�=����"�l��A+C�r3��7\£����2⽋4�$�xbUh$�{ۮ�����q^`���ōfa?Y����f�Y����~C>�k/��cq��1 N%Фj�u}���-��Vh*����t�Y��@���D�����%�3a+!��B{�,�Z�mdTLME���C����]�ArRRxN.��N%��m����6ró�H�r�O= W\Erz@�'�Q6�����z�Oi�$�#&�[�me�/���l0(H0�iO�>���(�z
,q�#��]z��bQ͕x���q��iV��4�X�:极ᒵ���"��X��ho|��g|?�Ԙ��~�"���Dy	����ťH�����%�q5|�?B�+�4d���yCh�ov��V�(0�Wb�ɵf���zlN�؉��"i,Op1y�ږ7��ܼh���/�H]�6xj�₩�.ۻ��[�TF��t��u�/���x0B�O׭?<q�k�S�2r�p����.�m���i�=���F��u
>�0�U�`!�P`�Z�[����k�ಎ����ݚhS��5�M�4������������8nQ���E���qW ӄ�@�̒��R��'w�:�`�J}K��2�i�Ɂmb������
��u�	���`N�����O+WpA.����6����S��D�t� �ND�O���=��Ԑ�F�2�|?Jk�SSm\w����O�]y|�t7�J���Y�sN�m��]hQ��&4p�ޗ��;��&@|�q3��'�x���Tm�pYI,���V-�?��R�˖��Dr����(^��X�Qrk������q���[�k@Ө��;'sm�#�|-�è�lKC���
��9�G����W̚���,غ�/\G��@�o���d2�vn�[��/��e�_�\q��ua�1.�,�X��wП�;	�guت��YS�E;J �m���0��f��Mt�VyL��7B��O7�����=�i�}GrQ�ϻ��D�T !�y�"�h]�^�YiDwF��S��0����z�T��A�R#���Nn�J�$�[I&T�M�H��>�h���Vw~Z�+��S�tY�nI\�~����њ�.��bKnqӢ 6���'I��:ɢ�0��>ɓ�*�;8�.//��ݩn���c�ӹ��-���N�ѿ___�"��kK.�Yq|��J	��	��WΟ{�Fg\���p�����!�2���ɠ�lG�YM$w+��g��XE��S%�;���}D�:���T�C��ի?��&�n��`�8w&����#�:>��I�PAk<��Z����It�O�����&���\-i}�5��
[7g*o�s��s8-�U�5����>@/��<:�{fY���Ƅ��,���L����"9;Jgˢ�ϴ*_5M���d�&��j�2�̇زYSx��H�5b����ǡ/�|>�I�I/j �;�ࡀ�GwT�U��Y���s]\w�*��}q�\�O��i�H�B��s��m)��q{St����P�_f�pC#E�^�  �ɡ�����u��VT��}d���m�v&�����@�~�*�����'N,M�UH�&�y�������F�}��?4� �S+��6{V�	��?�WF�(��m�&S4��Թ�\���g�xt���]����vV����ŔM� ��`�5��I�Y$ցf^b�j���Q�ߨC!=��w�5��H3y�o
�`�����+\2�����ׅe��K,w�xJu7g�O((9�1��.��B0��!	�F]��v[��z��Z�MtL�Q'6K5�E�>*I��=?��z��l�j���9��iO^�_�#�㤣`)�������u�Ur��,~��}�"�=
���l��"�/�~|�����~;]�K*[�S�;���$ʆ�́
>�
�e�8�&��!����|LNg��b�-�f�i�[}?=e�"=�!�<�j�XN��᥿���A�h�tz��gLT�,<�I8|tv����Hҫ�/ܭQj�����	ٰ߻P����@��r?C4��ʍ_�TM���]�{��ޗ\���?_�| ���3��N�t0��T�%v�b��AWlPO�����;|AXf?�2�|��S���{���C|�qL� ;Ff��M�U�B�xl��aW����|�
�*�S�Unh'`8�Nó�X )7�s�1��v':�4ꪉ�o���� ��d��Q��L�!Q+�5
�}�oDH��R'/Yf�_1BKM9�,a3*�?8���ME` 8
=�u��pϕ�#�|Qi�B-@}�|�� �g��m�H�n�/3�¹�ud6�_|�{�4Y;��?T.?|-į��4&�˴$?�j-RU����0]���B��+]��aݙ}5c�4  ��ū	��#�Ҩ1�i*�D�P�=�W� �3R����5]�@��3%��=��Q�a�7_MRI=�p�q�R�S��
�H"�"X9���f� 4�ɞ�vp�ˀ�N��o�ǆ�&��#`)$&j]-�<�킐�E��=o���7-�q_UC�{�Ͽ�K��Q5����',|rˢ<r�yD�e��>�Z��v���q?Z���s-���!��F���4v���8Ѓѳ�_Ϻ���9ൌ$��O�09�="U=}!�P��#	)&̯���9H���71�'rWX$��d!e��dyg�T�3��׶��AZ�̀�ud�y>ᗂx�i�9�_f�Z��m��	pN�-�5toڛn�H��H��nU����� �;�I����Z=���l~|�M�9��ۯ����p�����<?��:\�B�/4���<P�+ه0�χ��6��a�Թ󰰮1+��(����'$Un����61������<�t+]�T��mOV���3�e �q�U�N_��+Ch�y�áu�~t�Ix�S�
j�_��U��h"� )'�
�w�Fd`��&+����f��!�PG'� �]SZC�܌�� {SFeaC��ɖ��c�cfOM��TQބLt�J=�n�� HPp a��as�?�]�?�Z����P��bu�8��2�Cs��R����m�#~>B�Fc\����A
�us��D�NZ�y�%�8�}���REM9!k�:����1׆��[��᭑�S���**���ɖL	0�IR�zT��:~Q�x���������i����nA�w�|��Z�wHJ���v���Ө���*#	��l�0ߺG��򻐄#2�ItI�M�F�}�6�%���������cH�:�A��H��D#UR�R���|`KL+��&K��,�sMl��d���-tŎ�ꆨ&k+�����y�J׆-�X��ϗ־�]D!�pML�����%ݼ�[��ٖs[}��8я`����#�xc���ð؆5�\P��,?� ����4�E��+�ǐm�S����L�,�EB�2$��!s�"��^_M]�;��'�����[y���H�٩��.�E˙$q�n5x���~���A��*�[	��k�a����Cu/�%$��@��U�
��+P�r�;O8�����iV+���9OH�X�F�>#�aMrb/�ri��W1��Uv%	J��1�˕C�E���[�P��� ��J����@�@�kєXRC�so��g�-�������/����WQ͜v�pxz�@���~]��X�XѸk�y�Q�w�I
r}��e�3�h	��Ľ�L���-'�
�l;�QlOY�o`,�h�hf��=�Òhi�J���)��0���!`�X*!�.��4�6�~�%�g���t��XG�b3IK8��ai
���w���OTI�K�U&x���f�,�8G��p]U
,,~��S�$H<��E9�~s��Y�������7���A���k��<r��.]{����F� Gd_z�ӈ2�kV��@6���r���J�y�F�\4�!��Ǿ�JHQ}�<O�(�d�� 3��O�NN5==a��u��@ <!T}V+� +:k3�K$��Z��T�KFIֺ�`�5��6#�;�����e��$_b�­Zd��Cq�Ķ�g@�
��#g��K�t�}�,���dg������Sg�Ȉ�	긳��A��7�o����+9)��Є��w�T�rK :՜�g�?ܡg�$��w��ϓu\�	�ȳ-��Az�AIA}:�rJ��h�:Tp)2q��_^'2]@��*N���	"h2z,K=���b�=V�nDZ�>t�����ؒ�#�����}��Οn~���� ���9��b���s*]�@�{��ng%��U��;$��-@|��E/�ܧ�E��`(�>��c�����;}�[jQaSB�4���6L�v���|Ë*�;��q�vb��@�f��1/���Ś0K��Iaj�l&�QVR�63��H)z�
#�ܝ.�+fK���W����1�B:���S�PX�d�����:�x���#���������_2�:���5��D�MH�4�9C�_I-��0=��?R��f�0H����*k>0���r�7���'A����wtԟcE�4#M���(�t��>)��YG��eKg�0�½��	��-��$����T��?E�a�I���w([��]�ѯ9���4/S�IV$�a�>{K}��We8�.����Ψ5�p�5}�%#�:A�v��Tr�rt�r>Xԩ`�	��(mRXi^��DUQ뛖��Jl�H\��{k3T�x>��+��Kr���{ܥm 9^�G>:V�c�̑�p^�].������Fm�pv�rD&�}�h�n��K���X��ӓ&�a�T������� %��oa����t��������Im��\%�_oKĵ\oj<Pd�yS�6�̯�Q��*Xqd;o�g�
q�Hx���鷍�9�wΡb��4o2@	�+�`qߖ}=�C�[-�� �GI�1 g2�����Rh�?�rZ�"<���ڧ�Oj���~ס�ø��|��d~�٪D
qk�q�F`o�Ĉ��a�BeNx��z�>S+�/�ȯ�"�p8�~9|;�2�X{(�j���-Ǘ*�j ����)��
K���u�'К���==+`�ϛЩgBy�8k��#�A�4�1�%��c3��x�.)Q��HNoUesT���&������/I3�9��Yڹ����� �Ü-�/�C�%��mv�%0�!�Ͻ'��W���;z3m�g�P��@�GSa�~S�O4O�%�:���hw����Z��v0۽�1�
9Q�L�P~��Wjbd��K��q�M��p�j��)�h���$�d!cx�`������#�`6�P�f՞�0�}�F�nhO{ŷ�o���S�x8Q������*?Xc΄�g��8A��2��\"=Jw�=ل� _U�v�����_x�D���"҅�6#~�Kj8���d`lb��:���}��z����{��$O���(^��:ɾ�D*�9	0�؛�_fi8j�z|��z��ri�۳6���b��C�u�}%���6�����H>]K�GJ�J����� p��Ma0{�}&r�+N�'�?�~�39�8�-/k"�F��n��	�����M3��\�BZ٧����z���y:�ȹn'��i�8ʥ���9u�O(�P��
%;���6	��k�b�,��`��xSsNvi��1�O�
}Mƶb�S�r#	���|��m0��[>��ix�lԵJ���\I�!{]d0�\����RuQd��Пl�.��0���!�;����p���R�9��+���v.�������xԦ�>��w��7�ڀB�.Aم2E��(���ϟ�l����u�`g�,S��j��ЂN��h��-�^�#]Gj\��y!�_O0�J������/�\��
�:<��č/�t����I��î�1�nF�)�:Wm�v�R�LƮ�?�]��<KkӾ��g�9'p�8����w�z;~ϱ&�O�������������+xM��.�Dt����H6fxY�,J;$󽳏b1<2�P��lm"����m�D�Z#s������+�'�?�F��|��'��A�@	�K�Wל��x_"0����_�R��%i��B�5�qp���gv۹�-| ��:J�Meo��//Ǫ3�,l[�y�e��Aρ�g)R' �l�/,�}�
oEC�h�8%5H��Z�p .�^l����Bwr³x�8_�U�[������҉=�4��pI�� �,��W�<! $ܹA��N���!�����.�_�0�QL
�{$���Y�,W�q�a(�uC��2#������a<nV2��:q�����1�q��Up�HT5��u��z�C����x���F����Q��l㦁&�߫O���7��Ň{����zG0uPp���Y��2`��u
�3��h��2����%fEf|����m�-yf���ɌI\S�5Lk�,��X��b�Ė���1�A-֫Q�غs�ޥǽ������k�킾��F@HlC͓V�#d�ծʘ[J�b��͇�������t�KwC��S�ĩi�5�e�R|=�3�3ƿ��ZGܽ�5�����b�/>%۝��v�>*0��7 ���+���|)��*�>�9K�߬���@xn+D�ݦ��j��3��}�Zy�� v�0��N��*\��1F��.ZU�\��6(���.K�_ј��Z�k���)A)�p����u�W3���k#��'=z�a��>���'9��M4T)E#!q�s�,���4�*��C�n6,tΙg3���iE,��-GIu?Ds���;�^U�3@�*���`�H��~�Ƴ��y?:��@��tG���mv�T���Ĉ�;���0lj�����8�dۡ��|.ъVX���\�p{��ن(t���챮�S-�C��Xk$��ڔC"_+z+�J&\�g��1��gH�j~j�U嘞T�����V&�<�%�j�7���Ed��UG�oM^� �-x��c��әCL?_�d\K����nU��O�庞J���d��O�]&#�Z�#�~<���N�@-6f�d-�Ơ`K�+:��ֈ�j�R{����_>31���Os�3�&*�]�dM�����BM��a"���9˱��Ԫ�a_'����f�4rF�x�9�"~�o�d�n��:�4_�G���"x����)�)!�mx�V��-���r?��Tz��~���oS���'`��젇w��ιD�����t��?��SJ@n��,w[�nk�������}(����-NBxX6+���T�˫���e�0M8Bs�+�������G�с�����x�o�)7��Ѷ�X�h�5t`C�X¯`k�������Z�}j;�	%"|� %�3���l�JWQ�J�����v�zѷ:�rLJ�w?n������K�;2f-> �z��!�K�ϊ�h���w����b��_L.-�x�,*�z�����"�7͹h��o��#EYT�*�+�T#�7�Ҷ��<�g��V2AI�\P���[
ņ����b|7��ʈ��Sf����Bai��m b����ӓ�a7�2`a`���\�|AW�`�K�=@�YN4^�s�Mj��{���9�(�@�%�/~������צ*�h!�6�u]�>9�;�f�� s��a"�yE�)�A-ʽ���rX�����eYǡL�o��ʢT�/Q7_����lGdZ��3�G6/|oY�},v�~�w�ra$h0c\)e���r�)��n�Q��)��p4�ٹ��kb�Ȥ�Pv*�a�f�
����ڐƬ�#\�L糏����%� ���{�Gm�t��S ݖ8�|�z�ȳ���A�1V��&Ed,cF�p5�m�g.>��`�e�1Mi����Ş���K�Pū��{�����x�U$�O=�aU\)��Wp�O��7vH��u����v.c��µ�wo��~�(W
QA)�\�b=��P�N;�vV.=-��q:6��%ۭ?bc#2K��M���P D�IB���7;�䞦�o�;�<�]㎆PN�=�U���^|H��=�][}i.�����%�36;���	9PE�����[�x�TW��5��8�,�~3Xutȋ���W�zM�ʑL"�̆��L�>q1��	�>� ��֊�T9�{C���鐟��xP�(�=�Q*U*���ۯ7�+Ҧ/�J`� ��&\�����@��^>�M�}i3<{m&��<�$qb5挑b��{q���ȁ�H��'y�vE��X���~}m@�y�ΐaUkq�8O�Ք�����!����aA�[\�JC\��	&���!zPwa��:C�����B�B6;���*�|���@��5���Ǫ^<�XQ�𙂘؋������N����s���7�ez%�@?@�P��+ ���r�c<���^܇d$�8x��6�/�y��y�K;�T��,�:oZ�`+7Ez���4�P�e[��r{�}+�j�}�R7�p�d>�a�u�����oE& �4O��6�W�E���tˇ�#k�q�`�p�R@�<b^
]Ќqz��vA9� <?݆��+��O�!V9ZC'�UP�h�X8ۯ��G}X���l�| �ҏ�	0�\��-hX�q_S�ƭ��3�/K�7��M(`XIk袆�nͻ���'qɊ��]:T��Ho�n��w��iK�%�Q�ܳ�K!#�0��:(�e�ܨ	��I��=��`ʘO\s~"8BUѕ1��{�{P|}u�Qu��|r?�E6�`=$���H
{������
.G�{O��1�B$�X�8R8��*E�����I�Gq譁����* ta+���Ʌ I�#�U���-Dѽ7S�<n�#�2h�}�Dk�O�:/}J�JA�o.�d&��Z�߱K�fУ8Ԃ(ҔM$�y��3}�M�V���m	��[�݀����p�����lRv^(,ɩ�̲X�a:���3���DS���Z���ڜ-4�g��e���r6�CˏBsǧԇcf� ��k�Cm}��_I�tj��z�W$�Kܟ�L�ѯʫ7��dHĕG�]�K[���=�D�ǣ>P��V�0��{:�H�S1\��J��a�e�DP ��%|�I�uR+%=����U��`�L$1���NXK��@5�rv`�}T��Ǝ����r�ѿA���!t,4�vJf�U�����x����1x����NP"�6#�:�X�Y8�V������|��qPjl�T�M�KL�� ��u+C���}-J*A��n;�!�Ds���z�t:6�ɪ�d)S{z�x��Dhm�-�F�iU8<�ڑ)�6��U�Q�;����QZPł�\Qu����?�4��8h���D�p�&v�y�*�m�_t<<�G.�������F�~"v����>���#��1��QYhA�S>�v�P�>^C�v�2!��ԡ݂��c��3��lR�Ӏ|þ�� �!5<9XR���,%�[������0�M!L�u
��kd�g/�eTc_��z�Bk�ݒW`���\�W���-L8�>�ny5�(�>���뷝jo��`]}C>D����s�
	2�G�o��K���#國h˖�Lz/0W�.�������X�]��Y��i/S��^��	)�M��QK=튄��KH���?Dk��`����R4]f�ab�
h�Q�@���-��M�R
�Ǿ��64��C�R��^�*�7�޾�z��+g���� �5�����7���`�H�l�eZK��T� >�JPlo̡,K=���
�r1m��.u'�n%!O���/�{0"�&5N&��"��8tm���k�`� ����a`���?�i[~:U���qche����գ�����Lk��F��E��K��)��������ɼ�'�όC�~�N:߁ ��=7 [��}<���G\(���SU�*���w����'�uq�#|a�|�Ą���be�q�D�f�/b�L���y���.�O)��PTcם�W9M{m������ �[E�+C
���젤���-�G.�+���JC�WN8%p��1�.h���]W: E��1�<
�m�J`k�,�&|��H��&D�ʒ��.�Wy�Kz�bj.��n�Z0��#5�K^�㫳��f+Q4�L��z����m� �������m=�r�G:&V��^�l+
���0���*O���P�lbx�O&N������YpJ\��h��/s=(�����d�aF3�}'@iK����Q#������-¯U*Xϩ_`|%1sfp��ZL18���M�J���5(��z�����3d]�~��X<�%]Y��WWҪ%�d��i@C��el
����a��Ǣ�讀׮2���۩��X?gj�K��i�������LC;S	�7 "�S$�{��#1��-���p��y�ج!�C����s�����G��H��9�M�5K��-���u-��$ޯ_���`.����&�y|���1�K0�������=����TsBp��E������ibƅ�5Z�⡔8���K��Gҷ��������@b.Z�p�zc%C���U�Rw�@�u^�=��k1#����tפ\�d�
32�=��Re_˞A�Zp5wZ�?J���8�n�.H�]�̎���֛d�yp}��7��E�_Z�*vH@�M�5U7��(�^f�@$2�/F��r�\;J$����Y�j��Wz�q2�_};��~�8��zL�.���'Y~��s�h��v$�Dn���(����&��r����F`�/q����{Ui7W<�����x����
��J����@Y����S�p�#6�`�t�NrےW��Al8��1C��ȭ���4�L��9Bǡ�46�N�u��L���r�O�1�uP��t�Tȋ0�u�����U��?����w���^/��c���aj��m���@[p�4�q��/���IyJ�w�x�r	�G���ip}��{����1��ܡ�?���k�9sq��7�x�ΩҔ&!�@�Ю��6-��n�7^��M6�{�d�A�s�٣w�bc��r9��N�k��9�Q�ʦ�`*fZ����bʣ��Í��l᧏�=C+�$K����L��e��a+�꿸� �ҕ�-���������stc!��r��"BR��n3��аĨ�$x@�Ɖ+�<��4&�L�ϑ'+UH�~quɣm�n�R�dD�Z��!�jʣ�&~%�l��>�,"�',0)����Y5��L�/�.�$�}?����½B��1��t���,��^���6l���:+��28�	���g��x=��"A�������ю�,\]m	bؐ6�� �V����x[�%��.ϡ���� ���Ȟf`�����	�l�L�2 ǒ�W��P�fx�R��F"
�����եy�Z�r.3�j�y�EefS�uF�ʺb3� ����Q5��9*�]�������f��Y��"���_8Ļ��y��b��x�ͭ�����e8����!B!\1'��HH[�\��S�gӮʠAm�'J��]�nO�J�u�C����Q����"�ܺAHa�͞eF3I���l�-�U�=��2Hp�kO�"�>�w�U50ӻ����L��b����������� D'���wLE��B+��Ul����5���A�HOU�s����+���}��e�@�B4�7=R��y �Q�:�B�Z��4+�����tD�Ly�՘$���.C&�@R�"G<u���٩\}*$H=\�e���h�+AGh��ۛ^�#�R�7�FOz�LN�g26k��1ew�9G�Ut �4M�`�h�����W~�`S_��1�C 堯��ܔKKrY]��*=je�-���r&��$qu�H����t	�[Zl��c���]��hmӿ��j���r̲�e�3����߮��3�]�^�~Z�+iț�i}�WPEˈ�r�ٶ�3r���$�I����e� ��E�#��:�m#�o�{2�),�Q�n�H���F���01o�4v�M�6"�H]��H��X�g�Ԏآ\�'��f�e�U��S'�ڂ��.O�Fud���R�K��;7�J�}ѻ3�P����kʪ?�u���6%���〖�y�f��,WQ=��8攁٘���~W�P��������*�)>?Pj�ڤ]�`wā���T@��z�P8R�\^f\)�������|�]��gZq�o}dv������@����C�3.�c������OT{�/���Q�u��E}yj7����2�̱�c{��h��p ��{�῵�(n4'��3ۜD��'�/z@��d��:��R����C�H���hGa/���\0���,���%��<C�b˕�m���j�S�Ez�O�\�v�L�%���N��9mU��l-g�w�G:��wP<��M�6s�
�/Al�olE���Xմ-/�;X�u�lO���jx��Q�F�v�
O�����ӛ|�9"a� �9�P�(��o����?R`��y>�sr"Wx��}�c��H��SsK;S����b�*k4Y����Z����ƻ���m�w������,����E
F^w�f�1Ɲ��y��!��X��m�rF����Xr��e��	SpW�pa%�R������W�U�a?;�V9J���$�v��UF5�KL�\����^B���%!��
��5�D>���>����ϫn�cô	!��=}�j�Z���Cm�֏`5���eʋ{Ǫ��J�����2U^P�։�	��nv�"u���QP���֘��v��>�
?��̯؉Yz��Ǒ�zY�Ն����n��:K�oc&t��``0�)��&��e@~W&_�BھfONZ�F�!��y�6pd�+�pms��A\�lY^[��ov��D��G�?'� +��F�lT+&���v�X�1��ƽ1��ʗ}��]�I ,B J�ܰxX�cc�I\�]�-�uX�?�
�m͟C�������P�0ȲC-�@�VbfW���|�&X�bY���{���^8d*g)��<A<e�Ԉ�X�'1�Qo�I��E2��3ka����H����%o��b���*}㷣7ȫ�Xp��J�Q�s�a��۰T劅Ma���Ӊw�1�%=9tY/Ș*h��%��V?��t�z�}!��S�w?�e�贔<���(A��G��;xQ"������'K��H��L>��U�C���(��c3Qy0�Á�r�O~�]��NNJ��|��)���tq9�d��Bvd\�@�Rϐ���,��)�F}9���e������";5�iT�B�6����dp�O��_u:�d��LY7N�?&+��Q*���vq��_&6����in���:м��&c�#�cs�NR�����!,I�x����5嘈XD��X�#OӨ�\]�)�z��U��
��_JMI�"���W"� �~;�gm"E~�W�1���$��H�/z�r�Ǒ�����0@v'�Z�6�__d=	�������V��2۸��6 ��?ߕړg�.�u�侘��^�f<A-^��&���ш�H[�B��88}��3����� �Cj�	 K���h'��o��?�jJX��L�����|��?mb�MՑXп�P]�	�S�8�;@�C�Nw�4��YǇ9��Ɇ�!-R.i�. i�;��V��.>�&�_����/����p�,�M3��M�T��=B ��Eh�
���Q��.Zv�"ܸ��u(��;Y�Σ���4)�*m���Y\޳;�6Ys%���Q8�e�B�5����R���7b���MD�\'�#��
]a�xH�d��z����R
J��9]��쇌%ٛ}OY8F&�c���M/�1�.jJ�VA7[����kLf:I`��H�/z��G�~�_u!f��@�I9м�<���Z��8Y�Y��or��{���5��]��G��n1g���Sei��Nɚ�\�3e��7�]J�М�/�%�!�P�1��U�o�hK��E�T��94���?�4-*@w��[���xFab��Q�>M�b"��������/�t�ӟ4R�4H!�$��� �34^���?�"S0��~c����ΦЕ��7���ʂ��.j̞�$e���0ZZ���\!���b��3[L�Z<'ŭ+�PK�:�tR�մptpNgǎ��^`Ä5�0��^�6S�t���N&���G���P��Q��Ö2�OA����6:hIr�!��kj�s��͚bX�]��2�ab�o��:[%�W#����f���Y��-��w'�����3O;IKФ�揎�7�sՅl�� �C����9#.��ȝ��؞m3Cv2���D�ai�l�
��P?�k�)�̓a�z�TJ��X��L�̙�e�oJ[Z�bU&ᓟ�*FV�;_�C��b$�_T�z�E�"�7���A�̶��e�m@/
<�����Y@??97쉨�1�f�~�.��ηZ)gQ��h�h��8��x!��33����y����ȴI�[�䖫�t������t�f�=����-�Y�ýb	b��,�s|�UȽ���\x�2R�9/���y0���˘��s��s��5����SW��C~��k)l�\�(羵P*;t8��i�42�6�*K�\37�+�)g����8��V�?d�.�z\������Ǩ+T�i��Q3C�>/蜙w�b�賓Ȏ���Ʈ��y�+>CҴb�c{��T�^ø�����d]��=r���UHm�i|���R��+'hLU���9��~�c:�!���A^���>�8���۴?�I�h H�;��|�ǵ�Ån���6)�OK~ұp(y�+�v��O�T�!"����5��*;p�6�e�����z�8&	�b���Ȋ�#��픰8˺�K��
��KXg\����cT��8�j=���	���%	�C��w�y�&{��'�'p��c$w��&n�T�ɇ�\�Eƒ��#'���| XE���vjM���!CC֟��9��J|���vq��|oD�+�VR� #�@李l�/a��4|����N�7��1n��LP�qI]��3�`�e��*H�(�x�O�� �� 5�Q�ܓVu$����Y)�G�&x��;̕��O�;m���~ˍ%CѰ��L��q9�2�=�L혖�
r?��LB����ՆM��A� ����Џ�K��$p�8Y9;����m�U'�莐�|iж�
���]b�9�6S�%�4��u��f"�����+z��=L�;�hU8z&j�G�.��-B8����:�oP�mp�#�����!�+wV~];y�%#~�Y�l8�P,��1,�zߜ?齌CG��A���j׾}5���-�_�h#����6/���d�������:���:H.sD�ٔA0{%K�0�p�%�t1"̒���[a�������p�J� ���P���H��觏	������N�{�����`���ai�v.����K���i$�YK�W�ɉ��AT�B�����}S'�?Q�Vp\cY�}��,tbُ!�%���+��^_d?s�����<���?DΨ/(��j}�H��פ��а SXz~w��sL)s���j�09R)C�aG#����($N�U��s�j�������8r��a�ϋ����ك?7��)%b<>�G]8_�8`VmCJrm�D��0����$��$oay�vXOq����s�,s��NH%I.���s�E2R�g?�
|=����#���=�=�!�O� �������kblGݕ��Rg���v��|#w���^���}��E,^�[�.��*�vI����I��i	el��� ���?���4K"�����3�� %��Ϗ�B���4h���OS�^�Ǩ>?2@�iԀ%��Z �26�v�en�c�s��z$���w�ەq�i��+�	��.V{����,��C;��^��O��F��������ҋaಅ��	�6�� jUE�����@��h?���ǿ��2�ll�xql�:��o�R~�9id�j�nju�!��f
ࢊq,>���������%��bBz���r�o����@�w���X�P�CN���U@��3-�R���WJ���ӶP�y��CH&xGByU��IJ�.���%�l�oFɈ��ݛ4m@0���(��Z=�ş
V��G~���' �r�����R�G�D<Ƴ҇�U�.ߙ�@~�cXP��d�(�*Y�>�f����0K\Ub�D-.�;�_p!����;��:�&uʇe��Ϋ��nvQ\a�?b"��sh(ɸQ�G�tj��fޞ�Rb���xr4�E�r�^�M�lX2��C�i�GxГwK���~�
�kc��vu��0朖'=]�MI���H��'��x�u� RQ�n'�8��Z�Ev�����Tڈi)n�ܛ8�T�[�Um���pwvE�*6�Y_9���Z�y�?���Y��}��O�`/O���Ǩ�i�@��\��O�A��[!z�Y�yE�So��CĹZ�"o���׈��y�ϯ�|���RBGڡ�s,�9�*���[�@x�ո�V�׮}>{9_�6 ��mL�yI�����?�6sL���BSZ}���X����nH��ݽ��)<t]c�m�Aؾ��wq	,�����]��[saKً4�5�AS�l�{]���o.B�lV	�]���G	YǛo��W��yTGx:͵��vL�6��c��`{��ɨV;���*��^W�ýhaG(�M��"�m��%񯝩��Pw�>?���y:Ęi���&/<P��v+y@�������`}8$����J���ƪ9 >��C~��W�����#�mt,��I9�̚{�T��ˬ���[�ޅ�[���tm�{ր��v� G%�!g�!d�E�t����(+�HP0�V�6?Y�	֋?��tQ�gd"�Չ��)�7��v/ꯏ��qLs��eN�c�߲ƛ#&D
Q2��*������WG��p8�X֧ۢ"�c�M��#^�_�`Y���a�G�d��;;*F�}�T=�Yg�*���τq;� ,��]s
5S dU�1.?���*����EQ�e�z�9���v��2�0Q;����� �u<���O����[3zs]$���i�u�4vh�������h1�������_SWR�b<�ܛ^�hL?DuET���y��V���i�Z� ����)#Vk�|E�U+��iz�2$�,krn���#R���ZR�'���`f�<�D�)L���f���S���P�e�1Y����z^g�c���6�ZU�^Z���FP��mrM��������T�*�g�K��c�����=,���K;k�HFLaX�w_�,r�N��5���aj��<��Hۊ��f��$:)Rkp�C�ϯ���Pa�(@b�1���0P�/�6$ �hE��O����a/Qo�2�,f��t�ߡ0���u �����3)ѓ�]\�lb杖 ҙ��]m)ܼ�:��`e�-��Ogw�A`В�¼�^t���@1DR$}�^ע�񁖃�3�G��錬ZH�t�Eo%T��<�"�='�RC�{�pY	�a�w��n���.�-@�0碹�>;�b�������o��bx����aE��֬�Z��/��.P�yH�ͻ����ܤ$�w#�F�h�F�2��r�u77�9O��A����F�+�b���R�����b�l�\�����p��A��d��'��a��1*�	tP	�6��,׍���Jopjlݘ郲"^@�{.�E�S���G:�?���1o�*2�4~�	B�X�jЋC��`����W0e��/U���ilJ�[$W3�9+�O���!�Ɠj�W��4!��%"0�C�>xi�iXI�鼁�XhfziVXx\��I�-,�rvc���"��g/3-��7��'��_<�������o��Ok�O�ҙx =J�U �$�����/O;?�OǺ����^,���A�#���W���a�	\Ce���銛<��/�׻��XL��\A2rSG�s� �4��R�W�ZN�š�Q�eb�L����ߗG_\'�+�D\ ����.�H�:�<�]�F���%F���,O�J�#S2�uI��/���Fsg�Q��x���#3b_�Z#���\'e�.6�4�`��l���@�[p�E��B���ɶ|21�l������׉���4'��T��یY9F����C�O��k��@)?_{���Z�:|���P
/�s�n��!�@t�T�+��ȓcoSt��#`0Q��(_�En&�ɘ���j��8��?$"2�G�� K�(zv�u���k֚��jb^��\
DK�����`���@����N���fP/�?mѐ�U��ju߻z3\��4�V�82X��搒�?����$O�|r�/�|�x�C�wIP�A
7�D���{��l��MT^�xb�}C�P��Tm+l~S{�!.z�h;YX��S\Z\ݜ ��T;ʱ�~�:�*�E2���*�@��E����M�Pd	~��V�����J�$״�2�����;~@����UdHLl�]w�sNS_4���R����V�*�#�EcH�~�3�h�Ă��8K?���"���8OEm�}��f*�'�،׊�C���ځ�R�@#<l�\2�4c��8h��%���1�&��xX���M����Hps������u��Q�z��銲��E��A�3�0R�˂o<�e�?���s���R=���=�"y� m�U�^���͗�W��z��Ϗ4(PB�o��S.���9��2��kݩ㲍���Y*ш9Y�o\�1@o�l�C㢿����+��=*�R�D�����rl[<��6�`�����z��ȋR�_x�\Ͳ!M
!��9����ح �P����y��Q�ѡ�
S4̺���F�wʁ�8��UTd��%���N��i�Cqğ�;�r�˩���
��.H��K����7)�]�]�W_YϘ��J4�0߾V��Ӂ�S|�K'0�{_�Z%��@��^���E�ù�L&Ў�_AW!����3uR�Ӥ����e�2����1������I�Yw��!�9~ĝ���A[��I�����g�NNK;F�E�f4"��B�,]��{}�c]�6c(%��'���|��r&X.���M�Wq����$�w;�S�rH��r�@�@F��P��;�Ս���)�"�EPN�6)��@��i,����M�HSrّ>;v&b��}`�U�w!짱ФۜU��qׇk$�YŐ�������0s>��� ��ս�i�:�)+�;�ܱ�m(U�R(�3�l�� �o���6��	-D��X�x*}�E*,���	HN�t͢�kǏ0я)���>��54��B��AV���8R���K�suSi��ljV�&-r�w�/0������h�לPc��OSF�FU���Eᗢ[��^r�;%���e;��b 4��^	(��#Ԗor<�X������x���|ԓ�!�7^r�J���V��Cڥ$��IVE5���d��{�?�	;4���^g��0\��#I��] ��?���Y����Ԧe{��Sݨa'��+T��&�j�O���'>yߗ$Ky�1l^�8�\7#~9��?P���w�ĳ��&����ܢ� ��<C{|�L�/z��\ţA��Ws��3��fJV��L]������|�˃Ĳ!��;�,G�Bl�G�H�!
���[ڷ�t��>)���=Kd ��7()��X����l�[�-��t�ޝ���M�`�7����l��SV\�m��5�)�*>�6�p�L����\��aZ���0 �4��G���ì��>�I�T�3��S%��1&"�����8���Vd=©OfF��.�1�:�wO�;��:!/I�
a��W��{/��O�G�[�٤�n;�P?/yβ�^�;2�N��݆����k'ؤ�-L��],tʩ-7�r�.�g!�� w&��N���Ѵ\�hy��,�]�ͅ���z.�PQ�^C�!]H�=�4���g�����&T�0�qUY���l_��5��7DdO�o�tY�+�dP�qH�ʦCZ^���^��/��#��>�Z�;X��@{��KT>F8�FD���c2���㚓80Ҵ|�J�UL�o |�hIeB�źܝ4!;�&E��K��6��}sò��M ���Ax'<RH+��(�4�\f�=������4���	Y�.����R\{dU`�gX'�{��A�����,rC���&�'�a��
چ_����f6�!ps�/Qh(˔�Lr�d�h��	(��]m���!I�^.����=��D��S�l�O64��ۂ^7���F��p�`��ʩ5��6���+׸c����T��?)k�_ [�Ɋ&��c+W|��y��p�ъ� _��t�p����Dcޑ���.SR��oc�#�L�o�ZJU�F��:�������xseK�c��=�v��4S�_3�XU��#��Q��!�XDZ��lBJ{��^��q�^]N'�=�2��ތ��R�.�\����@�K(F��SQ*{�v�}�� ����SH�y��_�.8��5����;��#G^��%�u?3?xRx2t��?6�#��ƕ[/?�_�U����v�~�I��PMy�.�pޛp������<2l���hn5��X'�}�[�P7��ms��~}L�Q�q��D����仿l�foYk�ؠ��P�v<��'A)�r�H�3��;�W����}U*��*b�}o�B0Y�Jr?�)^Xy�4[Ȅ �5���I3��q�n;�sqf�Hf�L�}S¤���O*���6����|>�+��C6���P���؆D5�v�+ѯ�2���e||�l�����9Q�\@%���.R��0\��(�����i��`����yM�%����=D���A���׆�M��%)acd�+�H�D~��6�{�|�i�3����V��oFw��13Y��Y}O��׶~���4A�/I�J���Y�����u���M֐)�~ń����U�.��������@A���׻���(N��`�S���l��_���4"�(����v����V֧M�.�U%��:&$b��:�p����u@d�����	M&���1Z6"�m��(_��(=w
�)����U�ғ����q�"�����uj�Q�m!.��}�&j�_�����g�An �? �MC����F�%��YDF�>Z	L��P������V��\��Ã�����]=V�.�~�Z_�m!��W���>�-���������
��'�=��!R#J�K�_F�0'�ZǬ9נ���̵˴P�<�La�Kg���A�?�R�dg�U��M�)H@MX�b��.��%��Pq�����˂X�]"tȯ"�W�E���$ �K�ŰbG�#�E��O����@�v��5�ϻ�]X.�����=����?�2CMț��*
�c����"�|u�����
���7������6uqxsZi)G�d)l�LFA�mt|�/mr@��Ԡ��Ԝ0)��J��N�ʥ�\�J=T�����*w�� ��R�ey��V���>A2�^�=����KY4��v�bC�Z2&��S1�xھ�^jwnO�9�����j�LDb�t���S�6���:�/o����w�.ww��-i́���.�4�ռb��=
C*�t�oI���r 6�]���E_M�X2�r�}�8�AN����X��ْL��1w���?w|G�#`uW���MX���f����dEPl�!�?r�b9��3���TeB��A��2������h�q��r1��,�:"t�!����ku*N�Q�G�9��\
f���x�+2Rp�ک�|���t~fT:	(zАR��ߍ3J/��*EH$8�;_F* g�k���"(��4��:ʃ�0C��PG���������^�_w���|��B)�c�E8�'P'��a�ًBiV�^�lp� �ŷ��\߷��
���}�T�I=����pN�j�R:����BI�N$�y�r��/���%��\@��#@Sw��zF*�}M�a
�~6#�z Jթ���0('>��P��f�󊫚{E���-h�"�Ћ��[��k��+��=��S�~�j�$�L�2Wv�'��[���ϷB��!�$�Ja	*�5��B�Hq�Mo��}��������0p&L/�G���"Y�1X�;z��I���C6��p9�F����$!����<�SGm���f�����:������
>�m2�5� !4����k�PHKb�~��7�P���@��5��A�E1�E����)�ѻ��/g�v.K�οÞ' �em_��J�!��޷Tp�L�����4�Y��Ɨ�g�y�5H1�i�ˢ�Ϋ��<}����
�)2��DF�P^̽����{���ō�Lb�w �q\|�_q)$W�?I���9hV�T�4~����6H2�sqwX�0�}7��w�W�z��/1�v���8*��X���^�ѹ��c��A�͙�M�g�V��a��M^�y�O
S
�y5~�[~����k-�����������Q!E�}\�i*`�AQ톼�:Dn��<)	�`�ޅӅP��(�ۖRw�Jc:g�莮a�m����.��5ጳM��u��4�u2��lD����_>3��:~)�G����t�F�K:]q�H��>����;$E���雝Y*b��5�)�#�����7�Hޖ�0c^XP�O������OR�v�⹾<�V<�� ��.��F�4�BH��p��-��ʩ�0&�W���j�Ql�l[�r�Xն+!�I\t�C�z�s������� ���d�rhJZ��������x5W����Ѕw�"֫�/j�e7��{��J��:�������I�2�����XIX��f�5Dy��w��4��Y>:�jC#��TB����d�W���_:xb܀x:�5��8�?��t������|�Wt*^�Y ZG.��jL�6�jL���uu���a�����`�o��Sc�:���R� �[:���,卶������!6�C�?��C�_��ɭ�..sf��b��b8[E!W>��]'�@jY0��b
*�3�!�����.ɧ��7�[[�2u��)��Ct>Kh��+d;�����?v�	<���Ӂ�߉��[FRI��A�vh���R�V�		6?ct���Jҭ���N��OI^do&Fh�1�9��mT�M�d��}�z�pUX��Fu疐���q�k9mi�M��+e����J��g+�<i��	�Mâ����Lz���
$DJ�^Ħ5fҷ�ݺ�t��t2�5\�1p'l�+�fFt����'�I3YIl�p�(ϭ�Ü}c�{t( �sV�����/≮�*���V���@3٫�½����>���NiT�e��u�IgY�n��X�.��S���É�V�Y��jx`�^�%#��b��;�l�A`��&������A�������[$����6�);wB��'���g�]�C4�M���X�s�����H�����b��J��P��a��j�����T�$�T�A���U����w=� $����R�փ�ʸ���n��.���b�a�L&K&��jυ��e��S醘$���3p���H��8�\�r�_p�A3Nxr�x�!���F�^��iUm���ݛ�����OBi����c�s�����P�1H?7~o4`�>��o��;���M�s�k����?�c���Fq��]��7c�)O.��N�y+W@�Kl����W2��x�Fd�����`C�|aAS,k0*�Y�6b�q��ny)]!�mw3���I��v-�<�
����#�p" �������]�Uh[�?�TE�=��W񩫪2��);�Zd��!&m��jǍؕ\��E�s�N�jk�|�I��j#w�8��&�5� J�[}�]:�*���6T�E|]�s����:���X�Y�!N86Q��w\���:�W�W.����4�R q�U��B��8bc㿳,����t�d"o�M[�uٛ�Ơ3D�rw��bǔu{�~�.�d�r��o�I����Z�3/~�����a�����V�Uٽ�Y#��(��� 
�����l�!ͼJ4�D�Q���ɯB��ĳ,؉�:E��e��v�DJ�4g��������ߩ�DXK��O����wD����ԿϿP
�U�B��A���*�^s�
k��3N���-�ey@�<�h����5��m�}�����vs�4@�a(�S��j�+m�l;�v�F��������!�����@�+�)���BN�d��f3^)9f ��Ҽ������d�^�6!�@/���<���^�)l���%H��@$���F+T�Kn©4�Hx�6� �7E��D���8Lm��Y���Ֆ�Y���ql,��<� H�.���e�S~���b�&m��x�y�̜���CKR�P��""1Bp�����*�r>0�;p�ʃ5�SN޶�.�+������^�Eç̠}Y���2��������sӡ�.T���K]�yi�t���i�*ߖ*��Z�_��TWd��UjO�Pe_�N�)����T��YH�[���꽫�:A�ML#^��֑�u��.�t��So<�uH��B��V2�}P����+c�_��C2���WP�S�ş��*n�2\�c͢(dN:���;R����4��4Oz)���p��� �Zz�� �e���v�`��)Ì��R{��Q��!��t�`�9��M<��v�^e����}�����VG	�g?�i��+T�wT�$Դy�%�&S?r�M��Q!1�N����R0��6t|�Ӫ����Va7E��O3��=V`��2���9P?1?�{_q�`�f�,�5��T�R2WfVw�C*����J�����.6��&�F6F2���*��>�� �yߣ�acBF,C��u���-ZC�b+����V }y��e�JB��|��2�x�7�P#�8_�+�(�ؚ�#��h��T^�s��!9|5������i�8�k%կot����
ߒ�5\սɵ�7Q�Y���=�I>v�_�B7���-� OՅ��w���j���ʶ:FU5l��\�Gt�x7�*1�b?B�	v�ؘ���$�c=�lv;o��xC�l��E����i�B��*B\a4Y����S����9[L�t~Z&��E�����z��/
��MjޠT�Z�U6[6�����-����!��B��>�r�� x��59�v�݈ch���Պ���0�-<�X�
#C ���K+�'T�3�bK�ҵ��2���ϼҿ�4C��i����t�&�1v�8���&�	)��~��:�?m�A������S���7,ð��.G�yK����=�]�m�6��>�8(��}<���4�;�uy˷_��h.��(J�~�����J���_�'/��{�S"��IM���ዲʴ�������;0u"
��7PV:y��j�
����(-�Q�^����Z��J�|�f���@:��2��˲$�N&D�zKC.[a+�|��T{m��Kr~J��y�W��4��$26�Р�ઞ`S8Y?�l�)^a	��#�qɑ�������E�3(�đ�2�k*5F�ZE�9qUC�9�C&�RԇnU���X�����\�5k�&��Gmr�b��v6W�+�)U�l�,j2� ;���m��/� �R�j�����/�mX0��g]cm�������˼��$Q�NŪ��v��� �(�����$� ��",bp�kyU�J}`%N&��3Е��b�/Ci��>������Xc��N��(��8���ޖF�������:�p�6���`��p.Y�9q�IV�y�@�?�BSK�")��~9u\��@��5��č҅�S-l��p���s�\g79O�y��7�vv�	L�e�+�~��#�#cdfLJ{X�O��=9�)�xy�į�uQ��Eq��� �_O���k�B�,����tcd��E��U�"1D�K�X]f63vZQ�}�@�SP9�EH�`�s�c|1aՆ2��~+{�|�\bEZ~�#l���~��{b�p[n�P�֌��N�v���d��`4GVAN2��~(B�+>C
H��d�>��w��"�B�tz��!u���1\���&�4`Xv�����Qhrc�iR����q�ܟJ�f��!��S<��6��4��S(Y_B9���J�6��q��6�<92�}�&�駠�H����Q�B@Ȝ����}���r'HlZ���3� �
���fF	NhNs��f���d�o�,D{�<��,�Ȁ訢��rn3,�8�vEL`�
���)�-)�
P�`���8Q)�~��H�"�M?���+#�`�z�|3�o�q��4Б}@kVG@Iw+6ցK���mh;�v��Q����L)���k�|�W��C���#`ü�$�?�z���/��	����&�M �$ K:p�6e5%�,u@�+�&�j C��Z<�5��w����\����[�ɘ�e,ֽ���w_��K,T�fg�1X��������5�W:-ٍ
,��J�1�k9���a"���^6,�����q�GsDm� !�4Ĵ҅���"[���N)d����pNm&Ÿo~����D]�A����q+�1�/w9��Kb�u�K��%<��;S��W�&	��!�o#�HL���&�J��q[��Uӊ����Ք�P�p8}��焋O�u
�p2	�� ��-	�M�|�0@}]	���e��ys�)6ƱX�[���f�c�q1�'���9�+�&ky�N/��\ba䢮�V�~x����]�[�}��ǫaz��5����n@��%rJ,�Vvj'X���<qLB���wa`G�̂�WB�'�A����dfGƲ�7*���i N�8�7���dr��P��+�B^�L��ȡq�v��nfmY4`N�9��)�{M��CGT�o�h�^M�uK��)�G�RP$��Ƀ�'a��/�p0?���Ft̼�W�r�Lf��j���ġ�5`��v��.���#�`%��H
�P�"E�Bsq��SěY k��h��=��KW|V���4{��Ĩ�!�'{���w��E=ҩr�̚zm}=���%�8��rt�,Q㠢�M�]�%߳TL䀟syX�:�2B��;RMuO�ΩP��Z�9�~����i��M�c��Ԫ��a��.�^���ƿsNj�򔄧u�U��`���	3W��1��;ҨеX��! ��ָia��u�,R���nA=\�6%j�l[XT8�CgF��,9����w�ɻ��.�z5M$�WL(���19x���ݓ�OҨ��f*deO{�4�ϞKnWdEZ�%�โ��IXg�&��WԽ�K��o�g�f��-a�۶�VH�}�'3)�pJ,�d���ك)��{u�YJ�_��C�Z9��[�?�ĝ����ƒ.=1a��rn���^v�;y�CL��Ԣ��$�T���#�Py"�G��č��P��Kots]&ׄ�w���~�B�M���拯�9�i��NH���R�og'2���i���0r�v�I�KD�Z��G��b����ن?���~x\7��ƒ��L��"O��*������N@L7Qzv�*C@���n�?2)����>!�/��	��^�0lwt��]5ĭ�*�9͛�b~Ϝ�}�� �Е�����t�����m�	�f`q���,@ҩc�8]��,��V�7�{O�����"J*'��r�|��-�o���W��V�}JF�A��e�;�*e8)�K���dH��[(1<ʟ?��3�ZL|��y�%w.}C`B��l�\�_��Nϛ�R�*[7f�Г�u!䉒_?G��N$n��C�M�����a�F���s�L��g%��>>����r�+�%�sv���(=Q�� �D�����<�Πy�zC1���I��8���C?L��:'9��$����M-(l���(�F^u1��;fՏ�o !�Q�"LB�����F��y�^L1ĭ��j�x��z��Q�Ե�{e�0�rH��4T5��J�{r��؃9��A�����#Y���|}_����Y��?v��c���~��c@+Cz���qFVM)Q0*��$�e���K8m�R{�|�P���=ٱ��Qa�pP��\�^5U����`0!=�&�ik�����#�>2�vm�N�×��P06��O��2���i^6���ؕʻ���UR;;��ˉ
��o�@�k���F��\������]TA��q������ޙ2�>�%[�=#����@Ggq �9�i�{�'&�o&�DT}z��]I6����W0[pȄ�����`,��zhʁyf�+��80����,��%�Z������`�J��'7�]��]U������Rl%ė*�l����{I�Q�z�]����.����jA|���K�Y��N�~#�b�L��ռ=ϰ���� ���������YKl�L��=�_�-�~�j�IU~��7���F@�����R�G�~F� �b������H��QȌ��{;Y�?���ty���MZ��{Fx+�:�T�Jd�5�t�����*4�8JV�,Ip_�?��̀�W@|��ܸ!�h�%��z{A<��nLYʸz���p��5�qx4p�1�P�e쁼+ux|Gm�'�=l���P�1U�T8طcK,�-�n�9� Œ�AY�]�� �ġ��60�5F���8rXU{����
��a㘸z�ݒ3�p͓ZM����
{��#�
���.,��tHOk�c���gl���Oc��(~��ٳ5=����nXI�'C1|X�b0ze��4���6L���C=*Ԯ[��u9�d�.m�����V�+y��v�g�A��P3��|��b+���S[�%���:����X,M-�T�Ydl~:��,ᕼ�1�9ܟǸ=ܿ��ȇ��8m�4h�5  ���/�yƻ�`�\�e--c��p7��l�ߪ%S�c�cw[^�*Gc2`�c�C�?�'�ORbX��a�Y�J.�_b���w߽���^��>W�O}'�7R�v��u�"�/���u�@gA�s����hD�A��$�VlOGs_E\��,��X�@Nq���5�Z�9��2��N�JOl�7}A�1?f��b�������c]����T�{>X �M.��:&����o3�{�-��ƩS�X F
;��j��/�u?�N�㻛u��-S�p�AW �ѯ����B��u�ٳ�>[�+�vy4���ɘ7�<��/py�N�`��c(Y���i�V^��8�kR�ٽ�������F�s:�G>с�wS�4��=��i<� �XP�^��3�,^ȧ`�^��Q��|s��ejS����,�M"l��D;!餇��_1>�儂���fh�ኊ�O/n��Rӓ8F-�)�Km��;P���	'=�sP�
\�=��S�t��6m�������95���%1��H%%�s�F�8\�+�;�K�e�욃Ó4K�ɕvVb0���G���ů��pk=���6�^o�#4�?L̺,�柀�o�W���k��n�w;m�'fބb��=Ĕ��E�f��)�;̌�x�;.%\�i�b�\Q�_:�ΐ��X�R��
g����H`8�=�g�	%ҿ2���3��u���P`�(��H�¸�%`�Ρ`5VFu$g�c`�g�{����(n���Z٤��7�3�2����Z5�Y� !ų�~�^#�ƍu�9�/�BL���=�#o��r��=�܇�5*�
��S��0��YC88%��Y5]�v>\'�&!i���W1g�Zu��%����J�/i���w�_?~��M���?�5<20YyC��ZI���U���}BJf?��}�Zb3�k��^�R�輂���c�R�m�u��r���\��:ը�wSF煛�w�Ac�*̭#$0�N�~�1���Q� AlD	fh��l��D�\w���i>��#�;�������g�뢽@qЭ8�;hG��3�G%���JU9�b�D*�<��}i5\ȂW�L����	�ܽ���aǀ�y��w��yC��A�s�z�o�8
�����F 0VpY���~��Av�E�TyA��8��0�~���	\��6���#�4�޲���m����3tZ���������؝d�ltY�՘�'>���S��n~�I�Nq��-��Fv�>o���(�Kx�0�
I} ��V����c�ŋ��п7Ht4�6f+�����8�Y>���a	�a{f��Bࣂg+�q����=�ZȁD�f�y�ʒ���/��š�mh���xzӚ�_UZ��\���3m��O�+Ťهˀ�Zs�!����P�n�4�uU4d� q4�b���	U`���v��tEFy�D�]j1�ww	�g�s����}9?�U�?��4Ҿ�s:��D%�仸Rc�B��?ˣ7�y�\��]>m�s�)�jn:{��4[i�л�����j܀V�B���_�h�^��5 q�ܕ�s5��T�w��!����xK�y���d�ѱZ�k�"�<�|��1��H���N[q�h� ��:`�f�R�`~��¥�0j�2vt��6	5i.zpW�������sU������Z���K>&,� }�@F��K���1H�>��F���:D�������&M��v���K��(��ɔ'S���Ld6�Vd�����C5��׈�u�'T��ۜz'<n�bs�n_T
s0�xA���l�m�;N�T��ckㆾԞa�y���;�����q��� ���&�'��s�-nn�;�8��-j
�9��c@n�C��;/�W5hQ��G-�J(<��m{���N�-Z�,�V�?��6<͖��%�a*U�D$�����yx���o �h����a�^>�hT��d7�ǣ�q�@��D�iiu8g�_$�3�'j�.��)�*,�;Kl��O\���&��pcT������x���>'���ӓ���\���2�
 �ީ_�O#m�:�K���Y�����xc�7CDT�
p�$Ҟ���M���z���dD��,�Xg�1�	ö�>��9���+��XX6�D4��IE��q~�-��a��	��%��bL�y>�k8=9�$ב+���Z�i$Y�l����w�L�b��R��&Tn�H��9&h��T/�Gd��n�b#�{�5��n�x�e��z*Q�:��ezs���Ϡ	s�o��L<ν�Ca�۰Z���X?>\��Uc߁���C|�����Z��_e�nSpI�ڞ+�1\�!�jT�hW�i�$�Ե���-��#j��N[!lM�s�ʸ�m2D����3�s��n��ʸ�L
L�To!5�.�����n�w��eO�^�H�P���FF��d�@sO��y�����PT���cl�*����"k�������*�ӡ��%��9������<%��	������*�2�t��b�6Y�oo�%S�*���CU77Cn�+h�T��s�8v�晟>�{��5����]���8��.gZp�<wf��o]��D��H��y�~�V�*�^���;6��9I�&�A}-�;ٙ>��%Y��I���zl �����)ƪ��W�&
��BsY"_� �������&�y]�9ڮ�t���q����OKSm��-Pj���"�(TȬ#�bk�{	�ڬҌg�c>���7�0*=��Q%ܬ�5:t}�m��/���5ܸ_2���4��J�H�[�$gx�'M)��d^���	Xy���]��X�k�g��F��f�""|W��\���NPl��Yn����`/� ��Y\C��<�ͨ;HW�͕y�<{{�7?G�- ��Cdg�E�����_Os�t4�
~FNt\e���+~���护��	�Nd~nFU
<�b#M��	���U=1�$'��e�:��o�6O��Ί�3A��qMc�����o�3�`W����Cn���	_gk9�HE�(^#�T�eB΄��V���ٜe��&��w�W��K�)��[�B�ފJ���ʗ�1!
(�%�LH';)�h%�)��c��6�R ҹ�|�	Ti���BIf�0� ]��Y�o�Tg��C �9��=�Ҩ��}:"˝-/���8���x1͋��W1���A:{5�7�?�O���Ge q��Z�*'$�if{�?]'!����2?�tu�@50ǤvU[#�^�E<����M�4s(b�����J�<"�4�J�Ⱥ��*>��b�e�.g�� ���Y^�-��;�6�����#`#4�����G�DL��/���-��oos�Q^��&�`�-��/�^�{#�8��Q��7l��0����3g�h�Fg����V1�+�����e(	j����c,7�u;�eA{A�M�O�n���`b1�D���Ӿ��Aq%�@��Q���5�{�(/�P,Ҹ�Q\��w	�Y�CdHo��9lk��b�Re�0N~W>VN+�S���,<{?>$�I�O��̆1ҍ���2��/l�9,�Ɇ�v�
,�58k�_�9���>��qi��ϖ���2Ҿ�/ڠ�p�.�o�)񔽰}=(R:�	���V�خ�B�M����a:(�5�c��K"�������f�3M�50T��������
�GA6/s�ȢtVef�t��=����/Ww$*`�2)����f�S�.p*jBԜ�y�I�J�2�|<��RkB�Jse'uKk�y�PY9(~'��o�|��VO3iZ��R�x^��p�p���4T�̮�\��prH/�c�>!mGp"'Iq3��+W��$h����W��bRZR��6������|��i������{�a� �86������d`.�*�D�h�c����)h̗,b���zE���D�KD_nT7'�;:��ⅲ�)�CF �6� ፋ��A������n�QA8�z����K�n ̹�Ú�S�pY,��[%��_ܕOݍ���[1���*���S���Y��gI7��nQ"�
_II�K�q��)2Fu���ʿ�&���-�'��ȹ�x��,$�c�8r@�K�{=2�ee�L�kbF_����V*�/�"1�d�n��X�X>�O�R��֬Z�{54�j\�Гکr�8��b':�Ș��yȮg��AT�ǿ D&@KL������ �z�G�E%G����f3H(Æ�U��|���S�_!�8�ku��������܂��ft/��˕�$�}٨1�y� mfe��T���<W�z���d�w�Xd��y7���n��]K%NX������h�σT��ѿY����5���;�qJ�)�+�!���n�V+�O��/v\��%`#�d��폂�U>��c� ��$�	�ܬ�
C�_�c��T��]~��l^��&!���3=�*mGp����\��~�Bځ�dƑ!��W��f��zr���6�&a=�.�wX��iX��w��~��2����#R�z^a�D�؇��(�n������g��i�I��5���K��j3��E���'�C����:�<8��fo:Y�^7��h�k�73����`)�PBCĘ���B�ЇpH� ������vFXO�^�p�M
���I)��L�ERN��i��.� �j�~���V�hB�">L�dDMe��IJz�5Ԋ%DcZ�_O��Im~��O�@6�~�d��\ϷRR�������%��¬��p�ݐ�e7�����E���}h);���a��U�� �~i�3�_(K�.��pHu� \���y���l�MƳ�g���lL]Dˢ�c�&�XW���T����S���� B���fN����ro� p�v1�k�b���v��Fn�[i�WW��b���4] �y\�{��Sm#y;2LH��w�ɚ
�&5���L6��6* B_"6�Bv�C���?�[�a�j���[=~,K���d+��s-$\����x�	��Rŕ���샙�y���B](�Pd�~3�?�ccW#FY8�Zُ̹���%��`mn�R��mCV����i��`�u�~�����@�C�a��(��	7�����пK�<	�^[x�z������I;�������:G{!�bY�
*���O��T�1��W�Y��˧�A���Bh�X��ܟ�U���6��3�J��Q޲b��"�g��]�Yg׸6[ է@�P�M���`*����I�����CZfR�>>�t]����3��D���x� �̋���B>���4��g�ͺ����˘�XI������_z���E��aM�ةH���� ��M����l��O����x+X��dj<��h�jaW�=�y]25�v������o��A��GLL��E���[�T9����=���Xm��)8�!�* �O����&�NX���WK��#m��������W_^�K�e����l4ҨTDk ��1�s՟�!	�,⚏��܆���&s�dD��9�7��lX�RٷǷ2V;�g���8S�PN��6Y|�Zq���$�[
�zA��	Y7�1ށ:�hA�l�)�Ĭe�ވB\�=�o�p��$0Y�0����;���:a}����%��'�=C�h)���?�7�ځ�9��G#�QL;��+J�H���Jo�����E�u���'>�����}9޽��29���ҌL��/�yr3�~�DfM�%5pTv(����������F`���n2�e�y�u��b���n!���HI�Y[�^	~��~�t;�O)��v�D����������通P��N���XT�t�k�b�� M�Jн�G9d���l�n;��"�BH!y������rr�m�nW�56�7H˝�T�s_5��(}�6��h0�e����^��Uq����.��8���>k������K V��U����P[�_��0�<i���.��s��
���C^�6����C.�
��F/��׋����F�����rU#r�y�3��d��鯊0���y���uP��^�|g�d=T�bW������X�+m�˂h��2!�:e��G��th��"y܀�I)Z��ӱ��'D��f�\mb����R�굯U�S����![��l�!�-)vDwu��4�d7��Ѵ�~�b ��q���8n�Ԭ��g���\W��c%�8V���9Y��gO�,������I��_j�S����4"mBh�ӥ�
�􄊉C�Ye� ���O��Q'O#h�F�d���H
*ӛX�sU!�yE&=S�wc��@uh�r� Q8wEA�E��Y�d�T��砩m��&RAX �y$i�_��0��U���O�]B���8���ͻ��3�yJr��M� �d�1w�ϫ��=OS�_�칟�Y�D�v�����0���
�6�.Oȷ.��OĆ���m��Җ[W���6��0܀/��:��C��jb6���!�z{�
}�h��dŇ�q@&*ā�%0�-��Rl+��Z_�B�2�&%^ģ�`奐�%E�פI%t��c�eR�p�!n��G"I�S����g��?(SM�Npn��猂7\�?ˤbٍAqBAc1��ِ�x.��9��,��B�`�yb���'7�5�V��ՂX.�����5,GB�nA�W+AW��t��������ʚ��*9��e�QWҤ�ύ"���I�lܾ��,b~�H�2?<�-��sat�����vZ��������C~�Z����|na{P���>Ra Z�d��R�t+
�tA(^�X���E3VF����=.nX�php�k<����Q��L�ʹ���NW{���lL�`�����)��t26`��e��A-qA"�<F�S�Ä���1.z��C��ϱ�N�H�SQ��c�Dk6�*|T�uc�^��yw�3u+3@�y�|y�.��I_�P��m�۟����2��Jܴ� ĲD��*|B�y�a�!bB�p�@�vu��ɘ}%�a"j}Ns�yy#�X�EQԕ:�+f�8���n���7��:�N}�����
�4V�4yc����%0ɷtX.�u�#�./��)DJ��I���v�[ׅi����{Q)Gv����l}$�Np��1�T zس��;ܜB.pN�ɉ�;��e�<�@�Y�d��G�8�<�ҽt�*�䢂��/�a%�Sߒ�O(%Û�l��\�����T��MlU���|Ul��b;�<�-��3& W{Ct�+ >�>sb|i��3�_�Ug��p��S�JL>P	O�̋�]�L�ck��Y.hXd4�!q@lS.�i�6��:��al�yͤ��Y^����0��J�YTC0�j$P���.䥆Ќ_�}�"�8��o)�FX��]81�����e���:�i��TK��W=OkU[��*ΰ9@�`Z$�>�챈��ç��=���P��d�{����sҷ麠��h!!q;�����0pd�xz����}�)�ӣ_��-�9XV&�ƙZm2�5)o//�/��lMwn�4�ղUx?,�����K��b�s�G�i?�]��X�f�h����ƃ[���^���<{h��g������\��������7h�����U/�A�X�C�"\ˬ�OZ��A�F��J���ϧls�-���	'Ʉ�Y����|��˺��W��4<C~cgki�_�|P�H:�|�2�ڱ(֭~���ډ�V�`gR��� ���
���ivfg�ۄ�x�B��k��.k��1���_�z��y��,���A�W���X����u���;�=��řױ`j�'ƴ�~,�	�w7���
�i^��_`
���G��<�>N)�YF��@�` k��/�ŵ[N����&3�yr��I���/}��1+�4w����s&�g���Ju
\z��c�p��������J��I��Q,6hL< 3�).M���Q؁X6ʧ�>߳�'t���ix��1�6B��O���������X��/����)���ծ�NPD`��@E	�6{������E�١��H?�4�|?*� #���B�w-<��i	�-h߯����3l{��47��p;�,S�@C�,#��^��6���]�t�%��H�#\#o�9n��wV�B�\p�ڭ���pd��^��'�xq���%�d��YO��po@�Ў$<U�w�F�L\W�^!��ϋ�l����Z}�Pk|��]�d�Kl�i�hm�2K4��<D��P����2�itr�А&�<g7�v��G	z���=OD�&
�y����yW��M ���Z�e@��yԘ�����^,�~C��䔩�)q�j\�f[ �ҡ7�t��)����0�͞:��,���B)�
��8�EX~�	 .Ք����MS��a�<��|��V�+,N1��rb���J�_5n������~"�۪
<\z�L #U��)-�S�Zk늵� �w��]g��x�ug�o^{9��  �
z�J�Ln?Tf�焨5_I>D�\�J%��?xxׯQ�(��D8�
[�JP���NY¹���=ɛ|�t$��-)�Sp���7`�pa<����
(��^*�V�h#��jN�Ǩ���m�����JM��3���{6��a��	fE6��	"y��};�4JO�����̬v~�q� �0��L�N-��$�����AV�G��Tj2�1M�jE[&P]$��+<��ͺ曮]��b�M����qH�ڴY.�ᕉiD��l9�Z����vjfn%��|A�4������ŒFA�|�
���Ť�Z�IW�!�u�j�ò�K��J4����`?�� [G�������Q7���;�7�S��r~p�f���վڏN) j���[��Sj17��7��Ѿ���J䬨���)2�3�:y�P�mi�/6��a@�X�!���G�G��	�D�(��|����v��~�����5JʁO���Ć�{s&|tu��>JQHM���1�Qt ~���zF�ܰ�R���T!�A���!���tsF��)�emQ(�[�M{�E��l3+����Y>`X2-V9+���N�N���փ����_�Zt������u��i(ɇ��	J"L@eȎ�xZ�b#�X��=��2i�S�Y%V�r����D_s
�au w�d���K�A���#��KZ7��ϲ�\Z�~���3a�ϔj��/-��v�i;�Zq�~�1��������{���������:y�4�ϋ�
g�؝�v��+א1KY
�J2��t%�1��*�c�U�e�M�q�� 6�dy� vx��r�]�0��������Nl��ҕ�g
}Q��+�ks���	b(2���F�T�Ӣ�:���d�K�x:?r��I�������/�O��3\�W�����W4�T�XF�e���*����0���<=�+C�5�ܧ���9oU�S��Lܔ�*f��X	A���	z$�]���Sy��N�.���Y
��88m�	�;�J$�
CE���ڡ��7̹�;l�5�^�Y[l�+@d�af_CP{k��ۤ*V٬s{�+�A,Vv���%	���:�������rW)G&�z�܏�o��W�r�X3�Re�)qr؏ ����4�x��+�*V�:��]F��� 1!�fh?��~�[j\K�
s���0'*�"n�X����Ӧ�x��ԍށ=����5�a#0�U��\S:l�w-�f5�r o������XEpp�(�B+z��<D�5�
��*�o��V�+X�� �6��-�́.gm�?�B���*O٤7����}WR&�Ls���R���ݠХ$���ϼ�;y���*:���8�^1U/�J������Іl�/��Q��Ed��)s Ľ�W�eٻ�cVd?��}�I�)K��\I��3���?F 	��v�a��3v�[6�:��JѰ;-žF��������_Zv�/��%�+P��i�\� ��ʢ]T?���.�3$��(l�n�/�7B]���°�yҏ�$��)��I�)G���h��.��=0E�bA�"�O��߅I��W��͋�� �r������Ϙ��#/�譺|��@-�'��E���j��Aϲ}�8k��,͏/|<���w��Q���,$�aa����G�FW�?&�������|A���X6W��4�q�26�n�.�E��UZ��U��-�� ��\3��c�{\$'�>��gR�J�x 8��h8b���(�������/LH���I� ����^�yT{>���7����t�\˺Sb7Z:DFj*�D�N�x7�e����c;�J���t�-
�#��B�����t:K��D�0�W3-@�QZH.�	��ʣ8J��w��ڲ����/.��\�:�xR\f+I��2?�!�x�����Ȓ�J��EK}>��T���wѽ����ڦ�g�X$��&�Ti����|O7ޜm��V�8X$�W��������F�q_�=e>��rN���P1 t���Z�/-L.�RO��'��G�����Z!!H�Ǥ*yS\������K�*��v���5�Ȉec1<=��L]�1�Y� ��G��������n�&G����s�.Bh=d	�q�cb�U��:[H��H�iͬ=>�~�(��2�l��0���5^�]>F���b��\4
�=�!~$���p�>ձ��M8<ɇh}�6J�7�%��|(zϱ)8�tX�&�6�Nwlq��K����Scmma������W�|C�3|_���d��$KH�gN��e]n|���H�Wz(�����Ni>���e���x(NS��`���7��a`�E��W(eM���4��O�f8�]�dl%���%o������M�/��5��d�r�P�wʬS�w��і�h��OnS6�_l*G��4��+;o���dF�`�x�Mjb��"M�HE���Ff��`�#�S�"j�f�I>�߁��xy�w�?��%�Q�$pto��HV���&?{�~�	`�7"4 ����_`ډ��K�T��e��bJ����D�7h|�jF?E�_0Z������7sy�������x��fi��^ �Hz�
�����U�'|N���*�M<��9���n�l�H�:R���#N7:��8�tz,������&�K�ߊ��_J�ī�<(?�*�`_cz�z͗S��t&r�A�Y�:Y�:��Y��Ȗ� �5�S�SĻ�H��N���W;&��񹰋�a�ތ�|&��y�R�CHz4��[u����_�m�h�	�'��س'8%`���v�9QXA�9á�G�Ck�~G�y���)�Wlb6z���Mm�tn�K(��b ���������(���w�O(�������I���_bgN�q_j�<R�*�D�nм��߱�c�TH�=b�K/j>�a���[���j������=\�DOO�pƷJ��D{"b_:��-��M�/mt;S��6ƔH��?a���l���f���e�Kh�2}���z*7��:zbh?u�|n+=o6�B�T�N�X.�
�O��: �}��0�XS �X�)��7�8��!e���f90����a]��Y�SG""Z�P���(w��MH|1�x<�+B'�j���� 7�	w0�Ͷ�6��8���?n5aO�5fpn�B-��[i �ߧ�+��ի�]�L������m���j��M�{G�֙�1���h�Lõ�Hr+g]W�_2�0?H�u���9h�e`��Ѱ:Q��H�٪Z6�tr���뚨�r�S��'0F;e;�O���td����_���n�1��4��$��ݷ�C��`����ųJ���o}�׬WW��
\���'��i��tڥ�X�ՓiO��0�������@͠�r��3.xcͩD?!Ny<��<N	<��3Ӏ�����yc9+�a#��.$��Y�i�A>�c)?��#6A�"�4F�cM)�I,JxeF;�����ŽD��w����B�#W��G8�i�����O�Y��N<4����h����zB|�I����N5Qxˉ3#�4h�A0"��n[�(S�+�mG͔Q�1��44�G�����`��E�Jbf�;�ģm��Q����Ѯ<�_��j�_ŌA;��g�S�Wt"�n؊�x��x���� �� [�܄�7�>ӵD��㮦��C@o{q�g�Q�{�����\|,=��H*�m�};�Ax��i���]�=*3�r�"��Ɖ��vQ�$X0^��g+^<>�Z�j�����$�n�v�r����T��	Q���S����ċd����0I�<�Y���ՠ`��<��g����=׈n}ӥa&^�����,-!�j)k��(�H���hA J�_�G�#&��#���ф�/)��Kp)`�mW" �tIH{�P�\b��������Y5ֺ5�MY������m8&��?_&���]<_���?3u��p��Ĳ�My�`�7��w ߍ�g~,��S�Y�/N���w/�YR	#էݮ@(췻E��ߦEO2��m��	�.0-��Z���b���"A��Y�yd@�c�p$<O�6z��
�����1ϻ��;�ʭuօ�<~���0�� ��*��s��z�clͽ'�P���F���7����	.����n�Z%O�W�����B�ǤUDu]����`��$Ƃ��Td���\�%�)�����MD�V4�$�\��\٘�p�} �u�u����6�l/��	�L7È��ϫь<c�(���/^G�w�cM6�(��e]dI���:Hk�a�t��Rp%��s �c���
�x��8��~���ڏ�нn� �vJoN�h����a����) �?�������X�!\.\2�e��RA�+u��/Y�#:�$��8R�v�:�((QT�g>����	&�ѐ�eE��z���&ا�!A�)�S�ϴ�N��&�ǴJ4ȱ㬚�X(��gD��-r��잩���>`9���V!��#zOe	���mqTn]{78�_�K�9�t��[u��`V&��/L��\L�w;!e�k!��ج�8A��f�^�-��_p��Ó���t$�E��I�Ք]`�_�-��R��RH��A�~��mq��;� ��<�]�|m�eA"�F�u�o.jS���.�j�a� o�������H���g�w�a!��]M�k�"/���YuQ��+�"�}2`։�l��e��Mg���PvB�V��S�1qf� F���n�Z?F�lJ�\
-˘�fs%JZT�M
����:O��St��L�.�m�K[�	8�Dqv��>=�����$���fO�̶E����.����;7�����m�qw�\�'����:����5�̀��:4��' ��A��&x,l0���B;���s�2Zb$�Sen��Trx�;-�|��~D���s6������Ou�8$`���{up7#�B��'C�J*�[�r?D�b�R��aՅ�}���t�"��U/j�Ȧ�ʸ�;-p��[��O��ΎI*3�N!�&�8 �Z_�Bv,�����غ;����薍�"g!q�1ě�_)���� }XGScc�ڀG籥��w�Nҩ�a�!��.�?�4��H;iL��ܛm!�v)�T7e��M�Y�ӯ�ȃ\����J�Y/��A������d���=a��=+���8h��4��Ae�4�]Ԫ�WF�*O^ʞ��8XKDϛ���M��R��j�M
���=؅M"N�s]ڮ�<��Y��5霖v�S_��/}�	���Ζi���.O5�ƑMk�b�#86�x���VEǯP��/sp�>[�Q�ȣ_��N�/��勗L,�5�-��ؼI�~�^���х$tZ+��*����8%�o">Fx)�E�L�;��Km���*��1l�_ir<K����M�k5�c��6��f�Yi%n=8�p�YD>��͐)E��U�Dt��|�}ˋ-Y��r`Ѕ�9�Y7�s+w��9�����y.�'���%i*^2�F��i-�W	n��$uÁ3�d��7
x#�\D����ȟa+��!�%���H9�})C���Ó��\� ��K�B�xײwZLق���x�y�"��&����������6��UP��u\@{h��G_�4�Ʉ�:�μN�;pǜf �+����g�S�M���0؊�eV5!f�x�unm�f�R�R��cw��:�W)�6>.Z��݆�F*�y���R�me������GA�з̦r:f���竨�1�J�XY�/��Q�.K~w�Oۖ>�2R�ף~����-ͷ?a���	���av�xNƎ�ka¿ǚ5�F� URLL����ȭ��m����~���)�w����:�����_TR��c��i��f��a=8 ��
2�q�#m0b�=1?�����,�"mۏ���C�^�l���g��9�yM�|)�	)��T��O6	/NY�Md��n��j�t�\(lD�Ok����"�$?��Ã�v��"	���R�0��\��$�������?�g�� E3��k��X#"z �r��� %���>�ͮϳ�9;fv�y��/j�^E�����iK�65�ƨ��%Erl=?��AC�[P�B�$d��ɾ��'$��y�
�_ݩ�$�S~҃�6�Ζ�:��
?vB��iu�>Iw̜�J��ޝ#̳ӆ�(�RTh���)@:���j̹xr�jn��}�:]��p�z9J
{4��z�X�Q�K����=�������/	�s�if�$�5&/d��o��n��!�h��t�����`�a$n�Jw�u�ed	ok!W�3
%�<E�g����Դp�����cmްSAü_\Hoj�j�2�H��
��r毋����$W3d����R'�(>0/a}ga�J7H��nq�iB}Za!g�rPfN��]��ּ�����}Oh�1P��FM�E��!���ˏ%ݿ����ZII�_䮨!\�?5c/�=��&� p�*��v*hd�­���Ӱ.n��B|�Ȧ���j��8�)ܞ�aO��@̄����臤����P�'O�IP������t��I�(��)dԵ��j&+��(n 9���}�ܦ�ר/�Ͱ���y�ڄy�$ ��*��]�3�݊_,�n��ʴ��s��daJ�%�E�ߓ��G�E�sm��
x�Z�'�H��>�%��xE�D����2S+С�X��X��g�K�C�Jj��Kc�2t�J���6����7�`�x�H�[@�z���)Ij�x���F�\~�_p���w�����˜٨o="LN�a�ի��0�+��A��ӹ��Υ�!N-�����;
�Љ�ׯ}�aTD�W�C?�ea��uN��__�Z������6u�t���=4Tv9p;���.��Ǌ-��R�!�l���Y�L1��÷$;�����!��#�<�D�u/�v��<�^Ӹ����G|(QF"��Z9��l�䓋�tŲ4���oB�i?ӈ�49���1���D`Zm���;A��r�H����q~�|��K`�t�+��yy���u����ʉh�T��m��5 �X��f��jW��C�� P�W���8�@�A$�-�\�:���@'L�8�btn-ƽ��$:��JB��Q�����Sz�}�JЖc�6�Lx/,��4���y�"�@Sk<N�4j�G�A~��m㞰v��Rd����ZQ�����n1��n�,U�x�=TVS��Y?��t헦~$������+_���s��l)��J��qU�6�ML�I=X;&tP�U��7�;�d�i�Zo:���\��qe�����F)u�J�M�m�Z>���/Z��t���ʉP2M�����)�j=y�N�6�~ߓxpOȈ�pV}[��3�ik���1��m��9�?t(s�M!��k������3�@����CH���|ȶ�`N�'K�h���;�	��e�����Y��"Ȱ�oV ���u��QAX9K"����}���>��O���*Ʋ 2}1������&|h]z�4h�	�s��<֢R?�y�w�	�uA������Yo�r��:N�9R��wU�#~��ܞ���/�@��JC0��7����h�`>�yIH�Faf�<����`�S*W�)���]/C����x������ �Oܢ`�`[�ToR�H1����P�Y�E����r�����J���?�?p��
��q"���@�S��;EI�@i��x�`�ey&4����98&�˖�6e��rC��ۆ��5-��_��;���WM�-0E����؏�8���߰g�B��Ry���ތ�D�q�'��m8o�Yz�� �MC6T����pU<�����:�p�퀙d�Ծ2�;���s$�m����ȉ͞�n��[������l�ٽXl'j��6 ER��SV9,��R��X������y����s�צhd�1�j?���ѧ��W��5c�R5�h��� (�/m>w��_��?�[���8�Ͱ���4���61�vb��g1P���XL A���JZ.u�/��Őw�N^l-^ ㏪CB@��$�N���a��1�ri�[c�e��1T�����?�5%H�3�%,��<�"h8[�J]K�q���O#��i���y1�����P�?����Z��}�T;s^U�P��C�1YA� O�	L�MJ@��A�fۦ0�i+k:�{�u�F���Y{-�_��Ʈ�D��-�e��l�g�&A�\[s���-��ˤ�>����
�{�dq�8Ä6���/�����JΆ'G��~��؊�@8�����e��B6j��DTE��1�oX�n��n%�nKY��ĲH��䂹�v;��"-~{O.		n ���aFQWkD,/�:#Rb|��p.�ā�����R�$���+�*��1QMy�����00޻=��r��_ ��9��U���^A������랚�	���ٰ� �R��K���"��t��Jg� Ơ��YKGj�3,��&��� �����^(��{zS^��:���x��סּg��������T�;0����er蔵?���I�������H|��oI�b����A6���Of��i'�z�2�ќ�Ge$e�l����C�t�*�p�n�4�pj��" ��<��W1��Ы���l�z�,hA�Ŵ��;˂���$����2s��&�8�T<ԥ�7�$��_�1Phs3Lպ����_j�7�2��D𚱎L���ͧMavR�_��c���^W��F��}d�=����o��&0y�EC5�z�yX;�AW�j��{*+���*qodw���iQz�J驑����O���VdHZ5�xT��$e~y,6���#a�?�a�K����Iѓ��/��;��2��I���?��#��Q�N��s�ż��k}ds�	-���P�Ϳ�E"���g��q𗙸DiY��?Ԙ��>�l�o�gfJH�3��A��u�m���!��qu���GDN�	���7�Ntg���� 9\�=�T8݈��oa������B��Q��r7x(7F��
[�F�t�$㬭о����2�,��#ʨmD]�V�J�w�|&�L�8���K�(��[�]�n�L, �ɒ�։�9Jc�ޕLʢK��2LD~7�&�&��rǃ�xDz�oZr�>{�_���,���磱0C&'���3�����Ԏ��76uRtp2�x�T��߮!ó���79�3��;�J
)�-��Yk��q�S �("�/��i��	�]� @(�?��C_Cș�o����ƅ��@�ULw\p�+j�h4����7��pɄW���3N�¨��4�'��<��؍�06_g�-�:�Y3�23Wߍ�Ku߄��R�]o�t��r����x�&�����g</��qnǈ�TMm�9����I����ry����J�v8��@��TR�#�X��*]��]��x�dU��p�TI�8��6ƒ_`<��͓:y���A�m��)V"b<g]�L�-��~-�0�R�������r/���~cy��/^��噠�F��a��	_��dA��M��GBrKB���+1@>F���%/�����Z�Iǜr%;J�b8�Z1KU�|�f�P�Y�&L��A-�&��IiG���;Y�������>� _�0W�T��r#�zR"��ů|��8+O��i^��f��5b��k��k�"(-�)̯���&�� "%#6���5�{�mǋ½$�m,-��/�y��@{=�pD�����9�������!U.���������j�F���i���o�'�%�8ˈ�أyp"�C��_�n$~��J�z	�ה�wH�s1�O�@������@N��|�9��O�r�����
�J��Bꗉ�z�s�s���C�d+�������O�n;BX�]��b�D�I��Kzϔ��m�Z:����� � ���{���C�,ˬ�!�%I�U�a���꥖�>�w�ϗ����V{��㫾�7X�9I��e�lZ\u�PV�5��s^�1���kTN�}����a�^�:�$T����nwΑ�68�/H��i�[� �H�e��*M�D�Cە�ӽ[��Yy@G���V�����g#\�w^A���w�;y��eCd�P]C�wSI�b6f�!�Gb����	��8�idD�񩛱�y���<���N[ B��$[=J�
��j�f�V6�|�f��G������T`�#9���5r+|����J��@jܨ ~J�:�q�������J\S��o6�)��i���S�|%�}�x��R)�@ǔ���m������\�(k[���Q[�{�O����V����JA����'^�;Q�k��/��18���E2�U��-�?N��:$+&
X�$7؏�V���`U��õ�A%�a���L�!�Q��R�հ�^S�h^��3"i�{�q���"I��2�ڃ��d�)P��g��<g����ʢ��ܮ�Xlh2Q���"��V+a��OŽt*����U�p�l� ʗ�ښ��se�QwZ� EJ��*��nx�n�cr��='��e���S�Q#Ï�?�����M�ZCaw����	�!x. ��:v���e���p��clj�YzeR��v#��h���`m���o~#^<�N��e*�,��z�{�vU�$f"+v�����}n)եL�e3��B�����6��J�Cy��9���wSkV�ܪ7
��#��$�8,��"�R�+��؅�� �D|�����]�ኰ6T�d?-v4p��&�D�awl���*�ѱ���gcӯ��b��+j��)�Є���<������|�RP��\��:��tr���	�uF$l���#c�- ������x
�ziB̠�c��b�D���-r�i��2�Ǖ��c=$�3��w��W/����.�>�e��G�?��S���l��lA�0�,��|Pީ_
𔶷X�Bٲ �Pd
�uW"�g��S�j� >TQ���K�#����H��F ��h��=��B���]������f]L�*��H�F����j�Cz1��f����9�N�*ҝ6m�1Я��UE�d������m�÷���X�x�������,�����X*��I��M���SO2���	qPi��ȶ�͜v���U���]?]�y���bTc�'S���(ѕ-�q%�f�� \��'{��s��+�=�Ѽ�	k�X�e����5��B
��֫I��*��+���P��is��u�C�n�ħ�o����7u�7�u���W �F�-���ܐ�����de5��U�'~�
���l��&�6��w����}� $ �@8��MoS{���l@ W`❕�ͅK��/Y���>���NŦ�~�Ժ��t���EWA�4���~�!�?*f���UJeyJ�䶄B�3����|�3��^����"�^ ����G����9��e"��nL	��'�:j�q�r�f���7���&��:��DLH�t����kqĜ6��mlՆ��m!W��|�Ig��lpf��z�KУ������(���A`�)c]8r̡����P1���G��ܔ�5��sC*�l�X�KV���~�� ��2��ϫ�_- 5i$�� b�}1��;*�Zx�<E�_ �+@v�|s�.��a<T��;.��|�i��R��=�8�@�á�X0:I�T4&�Ӳ�M�:&;���Z�� XY�.q��GW���{G���K�x�"�j�L�0�}6\�] c������k����l�IY�O.S��c	��$+yl<j��������ws�����^f���X�����wQ\���U{��Ie%'�6o���O;W�u�A�:����(��B�=Ѯi ��v��	��$����4��f��L�(�Y�xx���6�;��;@���.q�ic���j�I���>֛��7'���D,�%'��@߱|�������ý���eY/h�={yBnT��^����ɩ�{ۆnծa�G��>#��sBƚ0׹\W+	��o��d�EA6KJxcOIt�i�
�����wM�훶�h���Vj�����^'�r��W��]�D����ǟt//�v��e-��}5qhL����9�>�{zkb��Q��E?�@nj3�Mv�
"�L_�!9�%s��!j�z�	�r�n#l��J��U��-��6�Dz����]4����˚�iO� $j��F�-�F�a*��.0�&/x��-{Y�,�MO%?��*�}�Us�l����Xx!��W�2C,k��u�(t��̘�E��������(��V���3��_�f2��g��ScX��������-���K��?�T���R�s�2֨-ú��V�4ɀ��;Y�1�q�S����X;h+b_�k��ڱ��YKwC�X��`�p�j�����tF<5���i3CS�αk�z�Y6��_��q֎��4MD����dx�[�N��=)P�_E�"]���G�	e]b�A&2�� �ߓ����<K��Gn��_�'��M���f�Nh�61<]�̓X�Y����nL�VG^S)�7��5 ��CEN.b�r�mG�G�4d��43܂�i.C0F�k��g�_)0�-���-���@�eh���F�/�x.C�Ŗ���Mo&�1E�_�*��Pn+:3�ޟZ|�D�0��m�d����N�41�>U�Ѝ����7���v��p<m�uX4�KpMڥNZd���:2�Nqԣ�:(��5�����N݄�0M�!���6�3�aF�� ��[S�[���2^���s�@�=V��#���!�����9��,j����Ρ˘�}��=�h/&���^��tgțB��`����	|w��`��@B$�Ѯ�s��l�D�	W��r�������4N���xh�jymB�1�4!l�'��;Y>^�W7�asJ�t�(��y  �vD��D�x`3~�aeG��!�vmQ�җ�	��wU�+A�a�_X�����I�T���x>p��ce;5�(�*�-2���y���V\G�v���fS�ٺƯf��GT�cY�J�[,�"����?G��Z��0{��Y�.3�DXO�76u���T^sM'�ַ�K!!N����>�]2Ǉ�� ��n]^P�/r+���z2�c�c�* q��D~��� �r7��Kz,�T&�|��@��B��D�nE�gaAfc���e(�uG��#��d�����n��ꣽ0���s���!��*�@t;�/A� ��?�!C�;2�i��$��<��m����z����Ί��
�A�꒰�B���.-`�=��=�Ny��y��z��x��������ݟ&�,��.{}ԥJ�.o��q�l�^4��\\����;�h���f=C;N/�I�#\��{�c��xB�h��H4󘋡zkGa�ƌ�	(]��
��QO�J����^�X+�q[5�LP�#��.a7�)��hgj������a�\*�u��O˅ج��\d?�#�_�*��r�FS1Tr��u�.�Sd��1g^{�R2)ט����J�J�7S����w;S�$�w�Y���s38������8�?�H�I,3�� $7 Y��tRGc!�5f�%��
��^n� }0{ʊٛ�ݚ"ć{�y�[�Dh��Ӟ��۫	���[�r���\TDݹ���V�]jD��z��	;�����x�)'���Og36���''S��L9ӯb���B������{�J����P����;v��~���~�)%G�
$��Y�g.�'�DL�m�����-t�׻�|��૫oW�#v0�z�2i�o$���p\��9�q>����M��%�J�M�9X@�V�`PO�؁"�CY�]�Qb�w����l�2� �ۣZ�x��6��W�X��6�
X�~j�s-����#�����o�S�>�[4�"+�!mm�\������o|P�z�G�)E5��\7����a�{��tup��Mz���F���3�fԧ�1��*��lZNq���ҍ�Y|y�M^>�I�Pc� �![��
I�}P�����A��P�j�Fo�uT����ܠ��I�hGe��ݚ����m��@)RFe�&��07MP$%����z��{���ͮq�_SQ��G�(0��1�]E�Fm����XՓor�ಜ��XR�I{6h�<���z'�]�Y�mi�� =g�_���S՟j
�rb���k�o{�|��R��B͏�����y�]�����u�<c���}���h|Ì*	~+w�7@*�AFBa����lC����Z��_89l��j�w�r���y�-kX!|�|s _�6Cx�v��϶Ȥ^N�E��ס�V��P��TV��8k��0zh��(�lM"P�L������@F�ޘ��H�#�B���~�w�\�<���&����[��Y�P=��t؅�Y��3V҂��N����,!��C=$&���N#I-f�2��2�f�}�Tx�$�Y� �iY)I��ۢ����ˈ�:�A���Z*�R�B�c��+�<������S��^�iY���;N�����I�����1x���BS�/�d���կ���2N��AY�#+�N����S�~��7z�[���H@L��!1��esh0�\U@�b�7b��T�z��ۘ�@�~���2�8{�t�_���L>�|�*�y�ךF��K�L��*�Kl佺{w�>K�g+�M���4����F�NOF}�R�/�I�}U�o��>|	���y}3�	J&�
�A�֣�V�}�B7EsQ<{<":�#�6ފp��ׁӅ�cRg ��ե�)_%#a84Pؘ�lUk��d��)�+V��Q��%�VW����vp��sJ���õ�S�4��i����jDq�$�Ig\�O%��e�8?hlA,PM�Sk����*����4�JY	xYt�ɡ]���$j+6	�>�'PG�o��1����A�����tD�_��7~�`ͯ��[�[���U/x(����k^u�&:�H!+��Ǌ���xg�3絥�'d���;�{�&O�E'e�I�KZ���d�J��_U6V+*)��sO!��f㍸p`~&Z@ X��@����S5.&�����P�'�Әq7��?Ⱅ��)��S[Ҳ�&k���f�,���{�S*�Y�4���~��Z�	�$j1"�{ŗoW�
^��9K2֮�j�(�ߒ�Z�e��[�-�(��-f�}D؛]��]ٽčx@@�i��:"1���Ӌx�k�S��(@�%�y�Rzrn�pqy!��|M����P{;��M~���$�'��~�+15��YH�k0�M ��]�"Kw����6��˒Q�"�jSk��M�r�ӡ��j6� 1N��!����1��7~`��*��%�e��dܕu?���	B��^�B<_I��4p2U�3G����:�a�(��{��E3^�
[h�*���	��}x�\~r�Z++�Ñ�Swj�A�Ef���oz�Y�e6��2�8	�>�G�üU6�s�(�?b$n6���7��ah��zw���Q�#��ށ��-�T����KNDk xI"��G�QW�]q�G���@��"	��0*�y#��\����6Ķ�OERK��ރ��+��BŴ�k%��*�mK
n�sO�o>T�	���4�&��+P�@��bi���IR����?�9�GS`b�>[+ݶϊ�9�"o��-�Dy^��3@�y?���B�t&��9w~��1�]��L_�0E���Ѐ�
��hYW��E6�
����!��W���{�����S77�������2�h�0OӴ�@�U>s�$&�� 0l���2���z�]�t@� ��}�^T��]��$)��r/YOC�R��� �zI�}�!l���΅a�JP+����:~��@��܃�$>%.�wMϜ��y����u�]P��_�i����i�Ɏf��;����H��8[�}�{���lT��,t6�e�5A�}���.�j�>(cΜ=�6�2��Hm����ۥ� ݕ�L�n~�ZN�QZC��ؙ����`r<P*�O4Rl�,�M우D������H�vp�z���e�s���>�������P��Z ��&_!���"��z�kn�Ҳ&����iZP�b���u4w�kY��I�T�	��ZZC�d�~t���lo
����DR攗��l)'{~���K"�gEGZLl 
�Q*�/;!��
_9,+Y{��9z��D����#ϬL�ͧ�H�K�s��R�J�[
TK����½3	uN7pZ~�tR��[o�̮Ⱦ�L}�=(�5�u=kT�c�t+�b<m�zUΨMϣ����Y{yر��y!Z�q������{�iu*��(�x3���z�Z��A+�>�΢ �\,�q��|trq�^�2��f�d��ބ�H��S� �W�lz�ԣ��2F��',k��1w��6���'{/A1�4���w�q�e��;��!y�)��<�`�&%u��5��?/?��OT/��)�)m��.A3�B�"8H��А
���}��Q6Yba�E�-;Y?�����}-K"U� i2��1����^��-�V�|n��Oh H*0Ar�G�z���-0B�:!���بNO�*P����~DF��7�E}�14S=�V�N�HW� �c�!KdJ��4��Xa��9�~��My�ي��#N�U��d��ĸ���7����!�>��CL� :T�KD���r��:����.��4�Sq�`����T�1���
\�vI��ex>hlވ�0|��Wk�R�7����н���K8�-�~{��s���@Mfi�~�+��J_����Ө�I�D�hNG��iM�����堍���6��F�i�Ϝ��\�)$Bؙ/.S6�Q�����
֭y�L���7GT������>�<و_P�v���Ǵ`�@���{�O��E||�R��]��[���5%c&)�o�5���=�5�� ��4�CU�)� ��"��o�J�+����QL���5�e-C���&9bP����L�c Gmb�};�.�-����"de�I�M���3d��'��(,ʵ#=���PO��	����=� Y���o�`����GC1{k���nEC�誛�O:��x�2�\S%�����~�t�0tj?<S]M�0�`�Z��1�>7�T���4{��j����2��uK {b�8�[I�)PI&č�d]���)�Uh�I�MJ�\�Ea�秧�f�9��8���L��Ԭ�ѦM�2E�}���a���uK9�c'��N��n7����+D=�Z�}��<!%Hơ��-���>�;��cu�4a����
5�s�3��LX��HW����U���y����U�,Y�t�5?������2^�y�U���B�)���n�{*��Tp�h�o�Q�R��&�C�IncL!'�[�S'��]����.�I�����?�����`����}��#M%f7�z�R%LǍwّ#{�چ3���/A��]]���=i��Y�?�|MM�@�!�u�<0� ���Q���#����A��aB'\Rh~Q�ӔEJ"�����z�&��jS�=�?����+'�@>�x	k�yY�_���q��xD���f};�,X!lp
�ɘ�sp%͋o
q��ݳ������P��TK j�_�7� ��p�f�A��͒�k�^�]+R�4Ǣ×	:6�)�����$�G����u�W��.�7k��ה�<�'�,�:蟘ӌ�@������z��ZI��OX�"��v	o��|��FF$,n�А�YR'dĂD�y2B�Sw5�,�LP:�¤p5�tpݝ�}��җ�,�Ne
U�F�È���T���݄���)��>t��9(��/ �'jé'���n���0�r����SB')��Pv�"Nf��k)���A���{��.���m���3�G�Ez��ss�V�"�.@]`-w�z ܞ��+�����1y�9R�����;����um�VG���uOO��n��
�a�����ച�ꗚ^���㖭 R�8��O��=��bw|5h%I쬂����}�X��x5����;�S�( i���zh��I^@�����VӦ�姝Y|M�o�C�~W-�jTY��ʓ���/.G�z��1{%�M���F3)l��C���0⑏H��%��R������p6���O�)1��T��W�t��RqG����*�MBq�L�s��TP.n�}k -�x�t [\v%Sj�˝
�o�2��l]y���v����Lx�GӇ�"��R����\V�ܤ��⬌]n)T�^R�&��Ǐ��f����ܞW�!%�������*HP&#�,j���>���:#6"o��2j��9�bJ��VX���C[�AG=t`(ZDn.N�l�D>���B��� m9)��MT���c�G/�P=����J�[�و�
��x��gu�9<{G_�?id����� )����I��AB�q4��/hK�4E�m�k���y�B��y�L�|}�c��P� ���j�L�DީS	p�v+j���<b���`��f\� ��e��%�`<�(�$$X���xM=�����c�2}��Z�7��|�b���f�j$�O>�Z�$�uX�i� �ܧƤoĻ�����R�U�T�����Th��M�-�E��?��3e;�,}6!b力E=?l�KF끲Y�wb��/_�	����x�d#���T�/�b�Y�x!�'A��-���{`�n�) �Ϊ�Д��T�_����Gn�"5��?�F����?m~����i�v��*��!μ
$�3k��,#F$S����.�/��IMަ�Ak�Gi��|�퍸�O�4��Θ$�(���I��3�ɲ4f�(���^\�@#�{z�d�J��Q[�!�4l�ٕ�&0��"״gF:�+���"����@s�9ϵК�y?9?)��\�&��:`1��M��\��+�r�̤���-O�&'�{���T�����A|~M�t�-HNľ�����\ 恡���w;�!�����p�4�y�'�BΣ��%��i������u5�X�D'�ET������
�"��ȇL:Jݟo�ɨ��w��GEs.��Fre�K�:J8�J�gdv�혀�i��tQ��X�Ep������E����4�u����N���yA�����x��_Cq��x�c�]�4�YmEo�����Z��\���Lw�MmTD��l\V����7Ux��$��NFw�L8���ɄT�p�J��.�REV�GsKd�VJ����u^إc��\o�)�AD��/��2�*����WI�00�j�;d�����{ӬWPl>���]�At8�9���H
[q$E�鑙�m�h����43�<c�Z�rKU8
��'�N�<��c����<P�bg��a���б�U!����S��`q�n�Q���7KK�%��mڋ�]��R#;p�W�c�#�Fhĵ�^0=jZ�DQ���5��s�wʻX�:\
3�Xg�?m��b���E�+'4[d׹*���5�����B����^�@��3oY%o��)����r�7=��G�U�X�u�e���R ����k�B��d�:�>{�|���y�1����?��EQ�vx������5g���8�P����ݘ�N��6뜜�h��ɀIș�?t.��9��N���D�����X�쎷���)�;�����D��cj�̄��A�U����[�����]#�����Nx 㪚pǘ�w�� ��&]�j�h�1ƚd�Sy�!�	`+$�E��L�u���I�(�7)<���].HrԿ�|!�GKTr	�+����YZ~h�{GF��I�J'�Ӄ�p˥W�ɔ�x����J>.럺&]t��FF�fh6qI�r+58~1D�3�v�v�Z����hT��m�ab�Q�E�ƚ�$�x��GnR���
�ހ��'�fVW�+�CGfK~p��%�0�a_<1v�\�c�xt7�gQ�!O�v��JT���I1af���xKk%�x8*�(k�Jv�s�/T��H�si��Р�=����ٌ��_�m�>�X�����G��_(x ���M-��DdY�����#�`��2���{l��ڞ���M`ǜԘw3���v���Q�P z�'`����\�%����WA!�ƈP��?! �䶵iV��UI����<I����0�X���5x����7�E&6���Q��p�t��5�IG�~���;Q[1���|�-2�r*�	u�^�Z�x���*k�k	��)4as_���^��3�ka�<
%�2;�t��&��BY�[C��O���9n&5Q�3����Ɵ�6��WM��eJ�v��᫥���I�8 �_�t�~�M���>��
���|JQ�����.Ӎ��ʇ|h�szhG����?��I���چ{ҁ��&X5M�xP��1������P�s^Zs�Oho� �]h�jW;B�&/X�L��8���<��)K�j�B9m����KU�
=����:����άLJ�2t��	�\DY�$���Nn2�?�R���Xǘ�����.�=ۃH<>��B����8pv����ho��Z �8�ιFR/��QXq����El����{�-)ۛ��&O��;az����Gk���+�.^"�Z���o�f�� �va���pUF1<�����'љ��d�&�[Β�k��?t�H�+U,�m�u ��֥w��r�UaYN���2u1�|��$��.��"\���'ZY�#D�����E��U׉l��;��<�Q�^g���1���u���7pnI_��*�|1q6�p�Z%��J����`_@����D���Yz�x;�v�ӯ� _��I�D�tZ]�mA��:r��(�CLK����`eIAS	႙��<F؜��s��.]F���{��c4�Ǫ-f������$�����SR��b�d�5�Hs����".��Q�.��[�J\�/#+/g��a	ё�a��w4f���Q�E�StE-gw�f�%Bd;RZ�S,;�+]��F_yd���R�+,z����@�̚�n��~�5��){�AV�T�z9��0,��I����dr[�e(���~��U #�%*��� �[�
@�,="g�
:"'>�T��˝��}E3�4����}?�� ��y��Ig��!}�!��y��u�{X�X
��*�:�zD��`�2� �&,x\��`���F<VX���	ux
k�
_�a-_Y�l�c�R�q�2X�b6+��;j'�QD��9�� ��fu�\.�pX�ۀת{]������T=�Ç�;���ڏ,Gi�T�@�)��i��Ï��&!iX^��S��,���@�U&��S�Yj&
�����;&x�w׎.�|y�Bj�����7��=���]�[��M]��������ߜ:-�K���J��� ^���.l�3��,^��ei�_����1EI�$��j$�C���vF�*pb����O dR�R���Yr�\���]��cUY#�HO��šSDAOh��Z�B��JaaM�to��J�� l�%Z��V3U�W0�״L~��r�W�0y�|+�B��u0q��3�Z�mu�_�[8Њ�S�%�y,��' n�c���D?�F\).��c�����샶׺�al�j��� o�.Z�e�=���D���ՠ��÷ٽ�[ H�0cT��y�;�b�XF���&[��1$r���?���"�l�8�Tt��Dɹ �G��mz0�]�<w\%����ʓ>%���P8��t����"��+{��ظ#��-f2v�is�	ˋY!
.��z��>Sv�W���B�r̆�}jИ����J���H ��il�{�ݜ]g����IY�~����O헅��Ӽ�K6�տ�W�,kl��b��dӅ�u��O&��(�3���f?X3V�+�W1L�>��një0�����?x�t��P �=y޾.�u��E��]�����I2a��s]�"_��ʪ�W0���'c&	�T���X��	t�q���9��ؘ�t�'�\ja�A�Ps�x�;�\\x����%��%�J����`q�.ft��H�y�qh�28I�m~������´���D��M��]�{6�dQ�)�̐/���f7�����a����j����	���-�
��&����Q�s�'i8I�L�L��)>;{R�[C�?�S-�<�~b����a���!�}i|�˭c�/���#z��"� �ؔHk�l'o�9B#��H���af�cg'�l�-������C*g8i��Y��L�-_�5J5��8����Ks��k� }A��!���Z�y�:�qz@�2P����Q�{�__o������l[o����)u�D��B7^.��Z�176
�b�su��p+M3D��g��-Q�z������Bê�V���6�_�cUgF�,�ǚ<�1>HЊPW\���#6Z��������GY���i�
W���H2�ؑ�\�gyK���Id�a����4��Z��m��B�}����L��D��Պ����N�+�3�Qp��}�+H��|���i��JM��yÞ��1i��:Ƽ�$!f;N���6�]O�(An�,Χm�܁g�(��b��H�t�mj8��S�:_�[�M֮��i[�k���^���-{T\�e�'���#R�6����O��a�B�6 J�� qr�q3�=��<���k�ts$�Bʣ�C�	���e[�+���Kq�����3lk�ڎJ�Џ�D�1�0#c��SA<�� r�=�˃R�����A`r�����]{`�$�ɿ��_'���giY����+]�C��U�Y�Up���~o&{Ҕs�2�g�}�H�]���"@�`@Y;�ct�q�/��������\$��j�kbt�A{�s9��}-9hN�x;��k@���ۣB	Q�G��zjtW��g�-�rt����]hE�CiЌ��	u���+���5��H�����!��8�y��q.+�^Y���9Y&�D�b� IcD��)#F�h'#	�z�+��>O�5B���8���<�Ֆ��jLjog1C��O��4�/ �jn�p���a�����>@Ü
R^����B�j�ߵ�BI��$/,l�t�#4<��\�t�l>�K/��^��H�v�m^�p�/�7��p��q��h�+9?�k=�X�#�V��X��{���p�A�������i���8��"�-�͠䈛���U��@U��Rev�6�k�%t���3��Z�k���Q� [��T<KL�ŵ4c��{2��5��ٵ_�E�/bEh9��	�{��M��Î�����m"J|��5C;+���Y!iZ	^}��������{����4+'v'�V�����o'�G��u�j�;L�"�;$�a��Ȳ����ξ��Wٰ�Uӧ�9ψ'��(K�L푦�$:�[�ˣ�	TU𐼸����1�L�0��V�[�a�A?]<�����z{yy�s�����n�X����H�vH���Wk��x�M���� �&���}$l�M��[/:Y���߳|���
���إ���S�����:CpeM?p�"�v��i�Ĺ����P=��s�(�� �	�wP�궸��tQ4��|Z�?.�#U�g���]�#~׀��/�|�!��[�ѝ��y*F0}Ct� P$?7�QX�R�@�"5t���/��s�P&�)�Ǎ<���"�=`M�X�Qu�?�k�y�lݫ3-�0s[�s�8^��r;���M�/hY��1ѭu�����X��pW�W�(� ^V�N�P��߼V�m'����@':�Q"���u9������� ˲��A��$L���4�29O�1�z){E�6I����W�����/���NH
�� ]qA�1b����17>����
�V�D�IU���yH`�-�����lW��2(R'^��y�ҷ�R6�W dG?`��@h(��3u�P\E��Ui�n�ʻ��g���0D
*�/�����;����Lskf� ��NҚF��W���ǧd"W}x�������)���x������:�n���,�@iG�
YO;�
��ZH8T]��j���h/��Ѱkw&�O֮L��*,�C���L����p]�5��>�� V�7�-{�h|  �&��d�E{ErpM��]3;�XC�3����K�]�G�!�+�q�r�M'���n��f�eA	~54���i�dU74x�!�J�È~Y�4�m˪f�ofΡ{�}|����&?
����#^S0RAd����H랲��r��_"Nw��p9u�l��`m��7�&~8�
�c�烴Q7���+��.���{���ty�&ܫ>ex�kM����N�z�)����K�M'��U�%�����a�%K�ٌC�<tUeK�T`�J���
��)?+��BX�F�0�\	qN4�|Ӟ�j��_^�د����@|��o�j�v^�4��qf�aD0�w�ξ������@���|�m��+�f�!B�"�ޢo.&���4o<!��X���Қ9�/�K���jw�3����DӒE���ʍ�0��:r�����4�JXW�Õ��K�ݗ��$��y_(f��F�=�{��q��j����uс\ �^9����à!+�E4�Jh��#*tN��|�,fs=7��<��ĝn0(aj�ѹͺae�ǭ�2��е��>"��_Cr���%�������cU���e:�M���Tk��J�dH����?*c���nf��"�'�s����.�L�D��0��̍�'u*G�|h������ȝ�W1"��U�>��% Qb����z%�����t�;;�_���[LJx�?T�*:=,��������8NHT���졩�n����.U�
8%"��3-�~w���,�������� S;��`����'r�oq;��L��Ͷ`����������o(� @�u/��(���;���pZ>�d�p* �kwZv���}����4R�>xhN|�y5��J��SLZ���zj|�Y���^I�$��<�}bS�SU�U7\/#���$Ϸ���	��J����#�ܜ��_�R)0�-�O�@بiY~�Y�ڏ��lY�\�1��^�����Ǿa��8���I}�aT�a�0Y׬¿#Y֋ޞ�V�T�JcJ�ۅu�c��������d�c���!{P0��d����lA
"��rd��>�L�Ht=�{�}k[��u5#�h��ÿ�I2J�]6��$��ε��֌��D����S��z`]��X����1$5O@�8�K�P�tE����9�8���Z�M��9=D�.y��?^o��u�i����W���UMw��[#�$���И_qʾ<Nt�8�� a���;^
��lc�ef�o�=����!c��9/9��3M	���Gy8�`��_m��l��R��n�͂�[��H�۶o�$�4AI��A]��l4P���ă�߉����9���#��o-̷;�c}כ�:���g
3t��EPedn�v4Cu+iO+4{�:�:�>��L�>1��ENn�H"��Rn>�u���X5A�?��,�?|�I�����V���m ��w�9 g����B�#`���vˎ`ƂV��pH =T�pc�)�o�f<Dr�H=��)�m�̰����(=�FK���kB|;�ܰe7���Ը�A���;�XUW���v�
>#��|㌩N�ܮ�8���� �w�:t�}UBC8�,.�L���rw|����׌X�R��[�J�~=�y�e?m�b��1T)=� ���3�\t����W��n�/Mf��n�}����q�Qi=9-���A^#n�s�y��
�;���|O��%l���ܬ�"�^C�FG��k ,��i0�':,;n#�����|�Z����	ܫ�
49�]�Q�
�:ɝ�3u�B�fhj���Z����9\m��D�\x^�+�T& l\�@M[K�֔N<�Z���ՙ�~:����&5� ��8�8�h 
�%/���;
�f��<�i��|��QN,�������O��)O�n�Zm[-0�5�L��v"��	�|H ��k�	�pe�ۍ$N�9N~+w�vG��
߼ǯ7�=7_W�V��@h��ѡ��U��V2�qn��S5*����Y���"������q����L��@�/9<U�HJ�?Nc	p�s�˜*<r���e���Q�e��MN�.��wݣ�ɱ"�v�L�skޘ�a�� r��>�v�A��&KN�s� � �V0uO��;_	��T�]=n)�GV/�O���sG�aL�>����IDD�+����a����֫:�+�,{��bE�ʗ{4h
���vj��*s҄�	�=��:ID���`�gG��0� ��TA:O����Uk2T�^��k�OVt�Nj�>�ea�޷R!��G9���|�x:y�/sMv�)�7%�9(	�~3�p�W����d#wCBP�-K�s&�+:���_�Fm�´�J���/�-�M�7my#����!�70$�Inq�nL�+?!�ߗ�$�ׅ��?;�AT�m��:��99�:1���{�����{.�8����UV�*Y�˴Cň>���Ckt�O�
�V!&�-`� )�>,Wĥ���d�������$��.{����ti�cصp 	��Q���定���Y=戎��֝�`�5y���9���b�YKg�H ��+��F�N��� �?U��`z�aẤ�׮I�M8D�#~öi.`vA��7��J5_�4/��{��1�����H�2<��!�f�i�Hx5.@��C]���ކ�8��D4��m�����.�X�]�����=L=��ն�=�=���-��6;Ǫ �ABǢ�D��yc�G@�P)7�r��vUY
_TH�c�]����k6*�B��1���ebc��.G�� @�%��:쵙���i�5�r"V�@�\�"J�֯���eFG��XJ���ֵA~1*�������l%KS�����%w/v��T�n�S�ȼ'��ms r�rӞ{�4:�_�
����x�4���	��>"�6�1�5��e� ��_��.�(h�%}�L���4\��ܢ���y�鑠���<�P"1�8=��u�&�?�T�~m��Mmڑ�r�ˀ���x �\M�~�֣��_���������_)�e�9N�[&�l��SX�w�����`�30��m�ԁ47�l��È�i4�U���V8��(�q�}ovҽ!��S@H����c���ʃ������:�@�ލ�A��H��x���z/Z�����2�>��6J(���1!�i�J�z�����a�q?���<�ˮg����C{�(��{rb	~�	r��kv�*X�Dv�*:�6u���K�J�´a9i9�(q��LA�I8�wP�xY]A'�����#o�b��b/�_{��=>����8��4;q�f���+Tί���~qQ[Da���6�y�puI���~O�P�d_8�t�Q��S�)��У8mL���yܗ>��ࡣ"�ضi>(z_�gx�`5��/�kAq���?ƙ)�f�S�;��ֈ���zQݢ�l��g.�����b�m���x` ����6n�Ai�t�d&�&p����&*��^�o��%n�ve��7rƾ�A��;:���!j��N�KڴYy������N˫b	7��|�YID�ŧ�f]Yk�KFf�yI���OS3n5��x/�AFk�m� ��4"�G5����O���U#�௥���Ê���V)�,]]k�аﰆ/2G�~+ٛ��.�r�O�g	=������x.�Z��%%�_V�z�	�DQ�W�M�3�����k��1zQ�g�V!�����W��϶���nx��IH�v^k�a?��-��ǣ��WhI�U3�Jr$���`r$���h����s��^�C�$�|��� i�J���r�5���y]��h�wcj3K�ٞl6ȝt�.��?��j�����u��k,YA�|��^��KNܱ6�] ¬v�+�~�n���/��K�s*m��4�h���$1��WSp�v(u�xF����p���|-A�E�ck�6D�"³|<m��g&`�83�l	l�Rd��l��#�K+N1�Ƴ:��L�ghgH��3z,'ir��G���]�0T��p�F^.�1�=φzD�F��lo�"��`#+��r��~�U.�G�~{�\��A1�OM��N���Z�� �ܑ)���3�����A��=hq�"�v�z�gYY6:�I��C�%��^�:��>x��a�u�F�KP�������&�Z4a���R�������	�)h0�F"
����}�ڂl�~LE��jl�6�M~6��z�:V�����m@��)0f
�]Ѹr���2�Vm��K!
A5����|�꬛�Z��Эr6���d�-(m���;w�^BP��[}��&J���L@��S�M 8���n>4��}���0�c�,p�����,��T�����w��~�)�`�Qc̊��v{=����b�	�����L:�? �����=!� ��q� �#W��S��%��q�6��<���6�"��!u�<�Z��E�.VFќqۃ�\���7m3k��5|cD���֧��b4��ff�r����渘s�P���d�p5}�p "���yRS���1��&m���P}ȶ[�޿�/�BQ��/{�N����a?}5�1FR�7_�Yv�p�i�Y>����d#ٻ���$� �[��'���!�uǅM���]��6�<�O�-_�����J�/֋sG��nyx rPS�v����=�M�foh��=�d�;��'��h6���W�S�N�w^�Ưڔ��P�Os��zy����Fg"N�K���%�n��)8�-�i{h��h�0kL�S/��}�xHejs*׏�R��ЃI�BՄ2�Y�]R��7�=�n��jL�K߫��r��C��?�7�8��*��5ᒍ��2tp�w��!~�G������7}�熲��穞dҁ�K:��B�2�OB����F���Urc-�P{��@czR�6�4^����ePߦh�9�md�GS�X)��s�{e!3t/�%L��
�+dÏ_��{W'�{.Ndb�)mM/r���Mh�g���L,��v$ڥk�pС�H�nUjtT������g��2$�Ɠ��0u.��?E�X ��y��M�}�O_aA�8�2t����Cd��mwN�zYN�>l7�$���
��#�M�{0��UA�4.�8?�k�j����	J-���°r�_e�ɬs<�k�R�m/�� �e-�;�p��ӯ|T֨����z��sl�\l��H��R+ln�7�Pm Ʈ7��L����o���+�Q緵K�ՌLE��;�M��v�=9�y&�իSuB����cD��چ�����hP�g���6DU>�Sӽ�w�m��x�/B��w�N��aڬP���m��=PzWz��**i���+k��3,�M.�'v�m��\��:6�`(���/��H.�	�<�kM��/�<���R=ҷoX�L��`ƻ ��4v��	-2���V��	�w��B�8�r?^l3#S�Ri8�^��!.���[�䍥J��e�
�|Y�S;OFho��3��Wbi�W����6j)I��Eq58ڮ���P|t/.0Y��5��c9��R���28w���܏���N�����U��c�����L�C�o���r,�s6.�I�z8�I�s�H�u ^����D;&��#���(�����ߢ�#�/dڒ��,4%V�=�����q�Ȥp��Ik-F�GA�H�OG)t'�o/hn��eA���h?�§�mА����
�O���\�;k$���&hZ��=&$��y�������y0�3����aù/��t�R�*�<9�v�����$��a��2��e%����VV�~��H�G�����t��vH<GA}�/ƻs8Jn��HM��ׇ���O�$t]Ƴ�cU�#q�f�9YD��1e���6j�m��hjN�0;��[@��q#���k�@\�\ߊ�֍׬���� ��ķǅ�;1���~,�J�=.�c��b��IBFĖ2�SEgS�@��};`	A2�����z	e#:����Sh��?g���x������p���a�{٭��+�P�W @tܣ���[�{�CI�h�����O�
��,��(����JVl<$�ԧ\wn�����+r���M�$�9�F�r�O8������ΥR���befl�䧯�E�MUzRMv�"���~�/0yE/���5k0���)A|��Q���c�?y�!?rs�m����"П8�ox7��ಡcc_�fLh�Eƶb�_�L�u�)Z'���LC+l�50=ug�d(]��|�#��H�0���B��R�u���>%������ϫ
�x�#��RCgI���}�Z^���ռ���
���)Yt�m�����-��6$|���r��a��R
{�*@�}�=�88�X&�gtK=b�
��0���)-37Қ:�!C����!��T��DN�8�q�!���R/��;�Q�����}x~�QSh҃���i���?�.�p��n��-�R�:C�;(�&��U/�.#�c�Y<�⇈�}3G��9b�[���� � +�_"�!��㑰���gU+(�(���xnD��k��"��t����(�޲7κd�xc�)���G���u*s#� ͝�~�C46Θ�B��LzcGt�r��x��6#�����m�H�J����M�q�p�C�&���<�O�g�����]j�E+AK����f�^�E�9�)t��ur�Ya�;�$g%{6���2K\S��V����[7/�w`P���[�;/~%�۟<po�V��A�q:��X�b��l�U���r��A��щ�	��7���~�P9Qf�*B����	d�P�Ap�z�ԑ<V�٬sݰl���x���StB���/�E�|T�m�T=f��oԂX��7�����.�m_ۆ�3L��.����s�gH�(��ǖR����4��˭N7e*�L�YS��i�\H�7BT�����y�L
xf*��7�gN����r�� ���-�ʶ��9Jn��������������zU־��>�1A,�ϧ��\V�����/����ۭ
h*� L�K
N�G�Β"l��j�'����������0�� �i�����0����µV�X��}�e)nk:�d\;p�MRID�񪵘s|�]��i���t�	�ct.(�t�~��_�D�ڟ�?������C� ģE�S�o��?��IL�6�*��'����
M��/mŪ��F�;�B��,�'��ޘ>2��>ce��-2ڃ/��}�ǜ�w�x����oKF�F>�����r㺻CE3���明H�]��"2���ZƑ!�+x�T��{�r.N�[�pu�u�El�{S��Q<Y��)�N�x~�%��O"��Tt�劔�.=iO�Y ���K��o�WjP�
q��rT�c^Bd# �9�:��yF��
����ox�C�A�>Q&l�����W����DDeS%g�uZ3b��K}�Q^�K�<�~��#�Z��%���읳�90�s�*�A|:
�S6�����d2T�2o�U�`����R��w� N�@cϫdk��Z)v,:��"��n�Y��y���"lm0�?�d&�kK���!|��ږ�H������cz����˜� d��k�VwI8� ��A�B���dߢ���c �?�K5������Sԡ�+#n�M�a�!|NֆŶ�k��[����ìQ[n�B�=����x�S{� 7Y��ʌ��Yd¼��JG�r-s*6Jg@@B��[��D��D��O�C��(.�t���t��WS�k�97"�n�$p��X�,� (�\(�c�̑�amp9�w�=w�cW{�b�]A1?�6���Y�o(1ģ�̈́nQ�Ք�o�+1,TV��꘢�W�r�!g����a���ٍQ>O/���k2l�2�6��f��Yd��u@4'�%d�"	L?��ZPE�3���S����-J��U]����� �O�]�Y-R:!3O�ln��}����?4v����8Me��[�;h+ի氬c�6k�ًӮ�o�s4�̒�5*S6�=H-֌��\?��o�fݹ���:�t#�.J��݅�G����^�Σ�f�>#�H��ZS���+L�g�����Z��*���G���.���y$���R�\��+Y�w�=\��(�P�9�&�*e���5�������������y��� z�� n������� ���G)��Hx�����u:�˹��R����@��*�B���Z�.��e:�d��� o}�K��D�E��=LO�!�x���c�\��<��m�
� r�b^£��7��q�U�pω�Q��g�U]x������"���R�����E�B�T�?����K����mD�.C��t(�-��<�}؄z����;��c!�̰���K_��S��:�Zvl��ԯ�,�wSټ&��X��Դ.�!i�]���m�:��K:��2�#��,;7E��H�����fX���H��gI�%9�8u�#P_A)�MY��� /�BʉT��l���@	v�՟嶕�45M�%.x'Ϣ̟�^U2n�quR=?ԛR�_%=�l��FҺ["�{	h�Ä�&�"�X�ߑ&N�(Z�����5�&�߆n[�ȖIx\A|Y�$�#�F�w���m��gg�I��z��5������Q���i�ד���;��fI�h1k۞.�r��Ob�(������>V�o�"��FL\��mK4��7������h�D�
���;��°ȐOEa� @�����2��P_ڷ�d��k@�y�G�*,�1n8U9v��N��8�Xg�)�*�7����~9�(�������Z`e4�������2�B�n�����S<	��}�#� q�k�H��7X��Vʼwda��u�(�2Kgx��ت)%'1_�vĆ]�O��.N�R��C d��Vϴ0��4up��S���N��_mT/�n��q�>����3��V���6�Y �3��җ��H�{�b/G�L5�Ϋ�c~�t�ɿ/�7�U���k�_�u���ZH�zԭ�A��Џ$ƅI/ �\���!�������	�&��F��Q|V��(�i/�<Db�G������z�����[���˻�n�r�����b�?��bh���,9^���	����8k�	�8=S/C���:D"��8&�V�2��A<�g����i�U��䇠{�#2+s���㦖���N����qGqMF̚���/�s~B޸V�S���(���5�)rl5t�.w���CewRm��m;3F���Ԏ�t
��ch�U�Q&�g$eDkm__z9�5��Z&>�C�g���=��ʹ�����%�u5{�a�$��B�S%��.
���t��FȚ�2F@U�߻z��6@ܫ�p�7G�]�e�V+��6R�0����&�@,#��hH�c�)b+�<�v��z�L�k��h|0|S��W��_M�� 1~�q<W����w�ΐߡtRaxAچ,_�����~g4�dr݋5`8	4b�pZ<���C��"����r{4oY$N��{�6=sږ6 ����wJ�H�Q�k%L���m�����iάZ̦3�l�-�6��O�ٕKs�R#v�����>fep�Ea��;;2�nC'w���F"�w�2j�nD
\� �-v��{��X��>��dWxP�buyy�=O�Z�� 23J,��12�)�y�����{eU�@8%��:|�~����Un�\��̓�с]�� ��K���Ī�37��-���)�`���f�σ��^#:�g5~�O+�o%���j��"ى��;�VS{��%��V��p�©n/�T�B�l�V����!�E;�r�w�!����#��vшL3�#�1Q�qqW�T������D5q��b���}d �\T�>�Q�@JEt��C)E^��Al�kSk�(�m|k E��paX�+�+�1���ܻ1Ʒ5���a�;����w�Å@����K����K��df��cs�"4;,=/�H��ɫ���E�Wx���e).� �,�6Hqa�M|X6S�A�˵�&��S��uDR��{�\�U\~6Ѽ���ʊD�L�F��c ���������{Yj�Ɋ6�Ͼ[!?QW���N��ľX�߉�r�,b�h���F��.`�m�x7�GW�%�D�ߗ��p�ȹ�,<)#�k; ���i9/��U������@��Y�O`V������m]�z!���
^,�V�`�SkV:YwP5fG�"��6����G�7:~��'j#� ���X�i��K.���?7�_u4�G�>��K��K��%X��(aиt�,��ォ�i�lFѺ���Of�vr���qC��gB`�Gfk�|���E���o8�q]��u�kxD���A����fZB2C��:W�Mi8(x�"E؂w�|ص���*�fT���a�^Ho�@ZA`����]�T�g�Ano`¾$�>��M��a`����� RR��*xD<�U�V�6�U5���^���U�&��7��*��E�%6���pK�Ј�9(�I� ��yZ�P�v
�D��R.�KU�k�5E��{��5	X]fG�j�/��6R��l�b쓥�gD�̓ٽ�Sp�gG���.I򏁆`�t%A<SeGI!���H� ���wjф95�rZ`G�kx�Ϥ�����X��x�>�3�>�G^��E�`��&�`�${,X�|*64� �O×��Y�.DWL�t�W�aԔ/��8&Ȋ�N_��=D(�u����=�0���K,���$>0���v�Z�we�ϖ�8{�-P��n4M,M�7��{��	�<��B�.$6K�P�����C�F���ժ�;0W7��}������]�J��e_�]�s�d�?�X��͹��a�Eŷ�;��C�e[ta��-��d�@�C��w�V��:��<��
�7���@�H�\����*��o�!\s��Y�$!��p��,�I~��-�����'0-��P*d�ˌF��;�+���:�'�jSL���f�q4��	U��p�K�o�ʴ鱖GB�>���z�����Ȅ��Vy�i��&�.�Fr�*³�b����"9�H��x���=W�}��	2��oA�E��a/��>��D�S�k�=��mE�~;�r�п�	i �)��1P2�<�-}\O٥��qmI�1i�0<ENF���q5�^S�F ǘ��t ��K�S@ݟsXW�d؉g��|���w1��qmLc���K��&��[B%|	yܗ��0u�L^E�uE���H2nrI7�?-0��H-�Du7:�Y��w����=&��ͱF"9I˴?&@k��m��ѭ	��)ُmPD�7��ɀ0����ٓ��~|!�x>��rzl�׽��+KI�z�y�0Y!�n�N�[��)yo.o�>7��ϰ=Y؃9�#��pg5���1��O"-�ě�C�ҍd��\9}*���@�L��bW�5�sf���4�ZVE����q�z����ثc��|M!Ej��@6@��i�W��RUVd��ᆤ��q���L�Y��i-�`ŭ�77�J�3ay�9���3^�s!s�f���$:��k
� i�1��|S�'q�\��a�,�E����}�O��`
�����.�_G4�%p���89���`J�I�F>�qrR���4qR�����&��Ȝ�,,���foL�T�%����C�MO�����82Yqc���4��O�tёm��Il�7H�������؊$�Ucf�k3���1�T�2ef�&�����l��DU�m��?��1>4�{��h/��
[���\����Ù;�Yu�l�y��ٗ�7���i���ZČ�+-��G4�u�3�+wL��]�����T%�9��[�!��~�������K�r?J��x��E����`��|:x�&F���|8	X�d�r1�8�/ٳ6oP�*�0��
S7~�����WF��%�2�W�����R�!�d�Gm}L�)r�>w�Ⰸ%h?RNU��9Hvs�Ќ�Uu����&W�Z��|���ث�p��'����+�
1���JcHm���RD[����4SeRn������N1�|Jlsol7 ����<���-u�5_��������of�O�eQ�)��7Ak|�����%�ʩ;(��U5�Y�ҫu���1&(R��i������<V���DS�0y45�w�����+��Tܣ���2>��5��ğ�� ���M�S	S��o���}�l"�/���!�!=�AP�cX �ϰ��z��Cs���($�{و1�O^g�U�j�e�-����y g�$���i�*ZoN�ԍ���˟� ���C<a�l���.$�j~��ݍC�������W���k��2�]|#^V.����6J��?�
��p�p w�ƾb ��V��_��{��ͭ�3�?�gٿ�H�s<]�E��֏��cM����6�t�=�:�W*B����s�����q��-6���\�ha�CI���ȋ��'"2��j5�Ҋe��b��E���ɳ�L1��GF�Y���A���\%m!�q,;����ώ,���s�7��t�5u�� �Y��.�W?�1L@S}��L��ި�H���`B �<ѫ���(cM����XĿ�»ǉf(�}P����\F+�Q���"�O������X�j�s-��o 4��Љ}^����؂��n)���K�#������NL�7��j��s�'��������W:��y�{�}�U��;ד5��v���	��I� ȡ�.���������'�RǸ��m_R���kk��n��_��a��Ci!�Ν�jf��l���N� �PӪx�r�]�f��!n�4@U�]�6�xw���F2vB�y�a��q�~H{,�zݗ�Y�ս��Ȃ��,����/�N#� lCȌr�����͈�M5r�����@�Y`�a�ѕn�\�(Zr�'4z�)��^�1�-���0�s��z����������7�Pڌ���m��hYA5��¼��@|i-��	���f駟�Y⛱2/���Lj�`j��Y 4)���)��~5�x����
Ӗ���1��N	�����h);>R������}Ͻ�O�'��?q��䔤KG��L��7@�%r�i��>V�-}��Ņ���ݠ|/k�Y����{�S-��g��AM+���tt?��C)��nib�M�/�����)"�RR���.��a�_���nD��.3s�>-*3�XG���:)&2Q��"��x���g ͓B����*jc�VLY��bIo^_��4�{8��l.�=�NQ��5\�N�yF<j�@'.S)=�b���})^�8*[��M6��~eF51�N+<fĎ���Z�s̍��w��Omլ{������E��(���f���cR�L��x�V|2K�W���-�ۆJk��!����6�x;������K�;5���5|���ۓ-;�]u��8u����&��XF?�F��c��ck����Wb0=_�ʈ���Z�S�uU����Pò-N�
P��Vl�E�p����`������O1̴�F���~~v(ƛ�K��gL���5�b}/�R~�O�Ś���B5�=ћ��F��j%A~�\�2�o*IX�j5}ʆ��<�	��P���,�|E�ȢW��ߥ����i�UKG!�0�F�0	i��a �9��
A�u"۷9���l�r��=��W�Y�P��}�o%�BF)�A~�S-�����ōǡt@aH$�ڸG��s��ꍻ�{:����ȃ����xn�zN�p�X�E�~R5�D��=�?A��SA,� �j�+�;�]��.P� ��&�R_��pY����������]�5;��@��M����f�	���ĳo9�8�L����kL�n��e�e�o�pu���J�S���-Z �hw7�p@���Roԑ2ʎ�:_�H�#MC�P��U`�z4|��4�h.J����4����X>�&�*ѫ�q�A��s���~AĿ܃؀�/������jDT5�>q�����C �8��<�P��'{>X�t��0HG֙X�B5/D�2�����e<���E)�6CL��{��^�����m0�o�h��_Ž���n���.3�+���eyGt�Y���gs��l,F0�4<t%��:��R�?�@j*L�|��	�ħ�U�(��d"��~ Q�h�UQ��86�����pe�v�>�<<�sm"+O����<@@��~S�1�3d���V�3�#�'������s 5C�A�M�Ϭ�&&ϗk������Z\�3p��D�v�V�1��Q7�Y6x��h�oh��M�5��*ʡ�F�Mݾ�I��1'��o3��Eʢ���O}uB���O�hp���2j�ɴ>�vR���Im����-�-f��p�?�^��]����^전LR��TF���1���9�H�DW��� {�ĭ�sWk	O9��D�<u�P�f���yk^������ӷ��+���h�G_~V��p��gA~+�$2|�VN�{9;+'N3~Q��D������>������6�a܁ :Jۨ׶K�M0����n��wWg��涮�2x�
 ѭ�G�������nAMo� �j%��� A�G"̳�G�Ԝ�����6�S6�b�`/���t��On�6�}���̚���1#�Y⾙���b�IxQ5�f��$����ē�P]C ��<��@��"�*�(;ӈ�W���e�Qn���6#B~��9����)�#��w4G�`�����t�
6�ꁾP��0О_?�F}�G&�,HUT-٧U^}�K��H|�ce��U`Z��#?�A�F4��'��+�Ń��S��OڈD��͸ޭ&�&�,-�p�M�u��F3�h����^���g!Mފ���kԦͨ��١K��[�����{���J2�Β��Ԑ��XQ��>ݼD0�K�[?�o��d	Un���SD_��&'����2�؄|���  �s�=�Ưk�?�n�y/;4\�m"�	�Hs�`	zLF���S�,�k�wM	�Mv`nI,�{H�fj�Z_T��o�k�i�d(���l�"a���>�qŽ+�aly�S�t,�89�#u����U����r��zx����a�A� �J�4��V��ᠴ����Q������>�x`��Y��fKttn��eZ����'4�'~�������~o/�tS��X�\REޕ���e�Mպ�(�r@��(��}$��c_�˙�XO�L�Ǫb:���'d4�m'�����N}wh�7{Gyev?�Ï^��Q����K�G�U?h�# �n^�IR�XY�ۿ����\��D{+5��1�L"S:���i'�^/�������YXLo�i��q�b���&D�ݐ���PX{����+*د�iܓ@�lW�|��g%�kdYeo��3���1�g����|��y!��Q��[4���T!��6�>�W	a@��Щ>�s(;���T��.�h&K�4xAh�ɷn]D��'X�N�b����&c%�W�m��R�z���X�*�ك�3C�.m�iP�v��VR�l��J�'H_wG�}rxJ�L�ҹ�,����M/)��csȵ��a���I�'�d����0�0�$����g�u��Jp/�6L��E�J�_�a*����͇AQ��z!���x��d���n}���u��P�@(rώ��O�Br|̘�x��:7�me2�}�S�?k2�,q�1Y\�<�,HK����5�hE��!+Owwl��<���� ��O�+�mA���v����&�Uy�~�%
�lT%�vܞ4z��Fg�iOy� �û��hڥT��J��j~�6������������q���΀^o�e�?��߸i��*%�$�Z�\�ҵV�ޟH�I؁�H����n!��"Q��!�`�TS§��ſ�u�����V':�a>�ũ��}o��M�A}�A
k�&TVw�F�J\�>�r���շ�G8
����`�����#�ax^����=zn�����k��%m+HV���~|󫚽3��W�e�i4g�A�V��#o�i�`�.�)��K��f�bĺʶ�7f��P�Zcc��uU2�.�$�� u�7�$)	��Q���L�2��aY�R�-be��-�����, wtO���͙�����������G��!��?!�
�kR��[�g���MI��	ۛ��G�1�U�v���$�����a� Ze�]�DȘo��{��C�y%�0����}ylj��ٛ(Kt-h>>���F����Lg�SAƦ;�6����#.�Ա�8��)2���?j�!�l�H�0�� ��vR��W�Q�x�6�$t���MB�[+��?jA��	Y���d�"�����bK�a��d����<ϱ�bxCz��a����l)����1��/�� (�e�+�!���,�q�!��Q$Y��0|�#�л�[�u"`:���ר���`K���y.�6��hNN"ñE�+\*r�A�}�-�j���'�b�x�t�qA^���R��|��_��8�@C��Ôʇg_��˅�̾;u��s��LW�j<-`?�l�Y�ꢝ�O��t�DI�;Va�����
:B^�����^;�f��q4[_8�����}�~eQ=��%´V��MEȣ�4�JҜJ9(:m�oȒ�jۜnpR�Ƿf�L� �(:���Ό�,^���fʵ��t��6�9��74��L"_yd>Dm����Q�閼��"{������=��e�h�5JWq�g��6��:�Ig�#}��>z�t�.�<2�@3���b�8�·T(����;����Tf#	6�IǻC]�چ�EE�Q(O�Z���JBU�'R��T�;��r�O�F<6I��<�ރ�:�G�Ӊ(-�����H�a}p�i x�:3@�d�f�k,�c"�ac�[��D_��1�V�tܪtE�F7e#����E����C.%!�_��z��`l�Ƽ��R {�����������C]����x즸y���]��#D�F�@Ű�7�iP����O���@+?�MRfb�b��k��b҄ ���wK���v<ӝ��,M��xc&�
��ٗ���O��1\��mAK�+��	"�.|�勎���r׮��!|���;��`���˺'#�N��)���?��!KO�7��^v|��7���_g�m��۟д'�0�����C�Nt:��M%H����Fc�d�.��<�)����w��'#��	��E\`��N��P� :��X"������C�^V[�e�c�������F�1+�'kk�)���U��LS�h{!S5�p`��?<�_�`����E��-fշ;���Z��jrhF�s����"�Tb��E��y>��:��R��"��A�z�a/��Xm�ٵ����2ঠͬ  iy��h/�I_N��$���!��ܻ~O�IH��Z�T�b�1� Y��cs1�ءh��^�cO����X�;�W�Y,h�(c�O�+L/rً���6C;�궓��'�8����ct�kcƆQ��c��6�	&;EB�IQ�P���#�����z�-�H)2�{��C�c��K۹��\�� �-	p����H���J�ǭH<�.�c���՜���@ɂG�m�V�� �/�[F��v�I�{������W>(�o��G�W���p���Z�N�B�*eJ�[\����h׀��C�f�c�[N����=��2߷n��`��v�pmR���0W ���цS��f��_<�he�����b�Z�k��Ԡ���?��;��T��*)ɞ�B�g�~yАm�ΈN4����Z-\����f�B�9�{�*Y�G�wy�ʯ����FJ»�Q���Q���Q�-�
z Q�N�^W*s8uz�u�E�����ίC�{��À	�Q_65� "��yҀ'Ie�������!RVx>,첐R~+4�6�W>���Cܱ�fsE	9
6��}0���Z�P����d�'������U!\�뷉��#f�m.w0�,���E{T��*`�Z=����4	Y�knF���W��B��4�o1���Z�r�ΐ(e;����P�_]��*E5�Ԉk��/��AWO5OLM�d���z��<�Nb���E>5�lw<P��K�/�p�YWc_ /:1�ݣ|�Q*���*���r�/�J�� �k$��Q@�8�Y��	o��,d�0�}�'�b'Ǝ��q��ɪi��)�i�z��8BJ�A�GӃ�a��!T��dp �#X���@��6�'@u5C*�y��H�T�o�Qķ��,���f�� ����YS��49%|�/���\#b����s$-�,���'��W�}W�[����2��gN�eٟ��G̰2����h�Z���shqQD��㣶�w��8咼s)�k�̤%#��7��8҃�e8/U�Є�Ҙ����Å%P���̿)���%���gg<���׌��1����C�?˹轭fj+::F~�2�|����g���`�Z����a�K�G9 |j�/��kg��m�;�������+�D�Q�/�Ѳ�-�Q�����H��:U�,��7����-�l�JL����yʙ������w�TH�,�}#�"�ARH��g��q1-o�f��5�]�J�e={a�#��P�յ5F	�.E����^� ,/�=+ a����������~`u�W���8uU��h��	<`��yw�:J_L曗T�"���;��W�j�nNL�(��i�K���n[�w��!�y �]�� ����
'�����TXk��0�ͳuĠ6~gp�b�E͌�Ǒj���)����fzQ��T��GǇXt7p!��c�,��۳�*�ck�6�ܗɴ��R�
���S���]
j�c���^��M.���T��O�7�1IWi��Eg�����T}���/��]N����./���L�_��ǖ���S��!e��G�R�����c�Ym�.�Low��'O�
����"�Ruϑz��?��Hh6!/�s}���uC�:ˏ���{���ռn�8Ƞ.-;Q���T��G����b����]�r	D���Q̮KgtDT��jk���\���Ȗ-��%Mn�ޝ�S�b{��ln$b�W�~pH�����w��ݲ���9�^��� ޘ��QC�tzZ��NC^p�;9��4E�VOQT =�;�P��5qJ�� ���5�}8�)(����%#!�GY�����OV�1�+�Y��B6���}d�G�Mh�� r����x} ;��_t�]�EC��~�9ܤ�?�ܬE�>)��-��.sG�q�Ψ�_S6hoI� �	۶?�u��2��w�K�ʢ�����
��a�	����3u;E^���jEf��N0�����=��B7�U���>%za#}�!���禉. �π����]�5zNC���?�E<���@�i��z�͍y�Q�ɤ��-��y]Ż�	\���v�6��y>�µ>��/x� c��LAU���8�!�q��c)�d��0�Jk�8���t� ���������>+���x�����լ�>��`Δ�D����t�j�a� ������T�\!�Y�˃�!�?��vQ�p8�Z��n ��*�9�Sl7�|��w|�M���VR�NlB���5,����=�}�`w!��#����3X��ǣl#�Css�U^���_z��R"�J�����(HO_�<Q(�].U5Q\��7cz��]�%`~W+�|#�m7dI�	JCh�`��ͭ7���Q����/T��P�Ժ����g�N�)L�Diۣ�L�=�v��i��AS��rF�Xi�lY5�]��j��m���<���A�w����/���7�A���~St�qc��Gh�^l�{��
�����-"@��h�=2� �%�A�V'1:������׌������ ��*`2����7�;���Ct�]��iJG�A1���}C1~�>�P�j���}�P�3��ُtV���'�|�9�"Ӝi��Cƹ�¦���ӕ>f��k��5�[�f�ƒ��%&1�λ<}�����w�HlQ������aHջ��02e������d] ʝ��9Z�J�2�u���d󳁜��dM��uf����jϡ�>20��+�L�`m�%�'���Z���2*D���q2V֔]��E��gCF��>�xP5�z�[iѫ�N�W{[�ӓ�6]4��J��ńC��V�É�BV���`���(7�.��=T6�b	�h�-k1��W���Gc��õ ��nF��0�X��d�Ye[/U�:l�x>����.��w�5Gx��'��\B7�BȊ�)G�q";$�Kc�2�ئ�]��,P�&�����U�ο:&A� [�"��v�se�X���n8���c�<��-ra{�+�h��R2�%ũ^�o1�2���j�5�;3I��r���XL_�9�ksl0��a7a��o[%)&d��g�bj!)�,f8�-��wDz�{�Y=|`ͯa,�8�T��B� ���5: �(	m�f�~�8�kcڹ|�b��ɔ�"
��P�����H�������ȕ�\��
��HFo�� ��&-�^~"���"A.ƺe�"�B������ݶ�6�QY�0Z�9s��KZ�9�sv���6�:�k�=<1�Y��7�Z�uʂ3���	��0i�L�<��,��
�nT[��ơ|H+G1����(�������	�Րr�������~��̕�F�v�g����uʋ������jh~Jl�?e��J�.�[��lNH�4�b��](�66f����,G���Qy��S�183<��k��G�b_JLMO�fj�4�%����^*Fi#�o�|��9�Ԧmh�����p��^�/Ɛ�@��/�YX1�p�-��`�buj��Ԉ=Ex���[�r�f-�y*�� ����1՞���e*�3�-�b'�	��qò������ݣ�7\��~�+j���[|{��9H�_4ŕ��0,%S�Y�61~H��p1�H�#W�(�&���5
���`7���VVӱ��p�#-wF�6��;A�l����`#7XtS�J
���m�%.]@�ǈ�6�]�s��gn]�X*��W�uc��$F<�\6�.@�:o��W�3�<UZju���$��2�q��H3Q0_H��[ҍ�;[�q��%��%J��XT���A����X5H\%	w�`Xȣ:���v"TG|�AP������ �R����F3�v���I�Z�QL�8>�Ǩ~CYV�+��&�9�5^s~E� �/�Qu���|>\3M{!H[��r�Y`�2�n�,��1���g���_A���5����Mi�@��,����#��+�eq}H6��1�]�P�QLi���~��܋��/ �,	MK��"��%��>��ɭF_�8��K�>Ö޴DKP�B4�=���
�d.TS��Dj������4�=p��D��n� T[+�Y���p��$�\P�>Ҁ*h[���!В����*���.B���K���Δ³�Z~F��[��^Z
mNo����QO�LF��A��Ei��ޔ�lv.j\(�T���(C�+�'���jB����U��^2j�4��z[�H�ACC8�8)h�n\aJ��O�=!��z�?����i�L�O+@Lk�/���&e���{�;�%1��\&��9*b@o��G4Up�S�%��)����A�m�^#��8�:\���HC�В����������!u|'a�T� ��>�#�6;���X��&�;������*�c�>u�3�e��g����4��PB���t�́c��;��u�b{[濕z�rӃL��/���Y���<4j
P)�S����\�11e�H��f���)��]���O�M�9���q^p��R|����U'<���;��q<��u�t��Q��j��ɧ�Y2��AY�}���{�٦�yB�e?[VW��(��ڰ�5�6�����aS�1�]1��^�}�#��Y��zΓ����w��0T�}���q<xAJ~"w�����z���C�����h���V��;5�-�����Z[�������4q����SWB������'M\���ܶS����ұ�g~���6(8�-j��?�/��(�*���]V�"Ev�F�M4 �5�%�
x�@60���f���^R����oA�{�5k�`9l��iA���",V�q��<��+�C@��	HjJwJ�p�n�RRux9�~s�^��}�W���'2ЧȊ>��� �C��a�{�ݐ˯�=)��Vqfn��-��U^_�M�
0l+"w���(�HZ>�v��A�Y�u�L�a)]{�N�����t���+d����f����?+�F�2��}��1��+&(6���evg��1O���4��*\�A]�x�g��?���9)t<�.Q�,�d����&n!λ<H���ȡM���AR�U���km�����;���Y�S� ���e�{T�J�*w���ֶ$�S� ��xʁ|�3�N9:����7̏�"�j���K�58=��:�uA���r�2CPw�*d���F��_<(C��')������.����ΡII��M�8TFӈ��a Ì�߷��uz�>E-;�c \ٹu@����Ȟhl�6����c�I��!�°��K�J��N���B?�L{�Y��%�/D�C_;�n����" ��Ѝ���V�G��zK!`�&g����|��mz���P�����A3�as\Ar�_�a�³��$3�W˪���j���l�����R�-��������2�^��M��[[L�o�̰�\Pt~���"ٛJ�Y��N�	��<��i��ɰ�j�%�tڦ�O|�'�:�9B��o���Gkyn��Ջ5M�'�:T��	w�$奁�s��t�Lu�,� �օR���&�9��$	:~w������.��TZ�Q�te�k1��o��ҵ�*��d��񠶸��y�r�/�M�h$��+����%P��YѷIT�N�r{#�x�G���]� �R��}����G=62���O��i��
v��� \^PP���6�j =�t�f"/M�˘�e�.�9�e�:�+5���Y]a��S���f���A�L�����I�^�3tl�X�a�)�P\@���
P���rN���^��Y�y�"25Z[o�ԉ��<��@��,>q,b�$�Ipk�>i��>>��NK��&*p�q���A�}�X(�V����f
U�>i�R\�\_4�)܀����J��f ti���=M�a1�2�i�˝�*e�������ds��C���a����/!�Ǥ��ڼ�R����\����_���UN��@9���
{q�Ff�V(��c$0����'��x_��"���~)�����6�$篐���eD�f�{q�=冬��:,��Q«�����di6R5[Ua(T��O��k5[D�rD���C?�����h��_C����qY�01�,tV7�S{T�\�;cW�I�;*�_��:/wJ���)�Փa�zynݝV��
�M�e�l?�y�?�&���K�a�VrZ{⥋ �_lD8�2x?ʇ�r�'��X�(��7�
@�;�HLp敵�L�/ȅ��u�&��T�J�vZ /!b���)+��;���wQh�5өyZ�S���|6g����NE㾅g��}�B+�u�,,o޷�R[�l�V�s����; �Æ���;��E�[m^�����~�MXg��բ�"Ȕ�#DaW��^�+�8T2#.�8�i��J/���
J���u%\���GC��#��+�>����ꪤXYwp:�$Cx�ۊf��Wz�DPK���fpO���Qj��v5�ܖ����O�Bz���kA/��n�9��HW_`U�����sE���GۊS�O��[���|�%�o�aX*TP��h��wM�ԗTҒ�뉎,���_��
ͅ��7�$@�EA$y>ET5B�tL��ln���\�#�0��ၫޗ�C�T �E�C~<���ٍ�lJ���#>LH�����ъ�f�^�Db/�5�/~�7l#dI��&u�'f��Wa(�d��îp:�%(�d��Q��-w���*py���.~I>¡�0ȍ4.Gz���߁:,�N]X��A@�:f�q����TxNw�"�,g��^퀑���O�*~g�"���ǯ�2l��vUT6P�V��0&ў�+OX :�����*��p�����. rf�#���k�4�8�,2Ur����NV��˂a�|�|d�6eZ ���W����\��2Pt�8�T�+�[�Sse���9g��K�PT�l��-ߓ��Ou�c�$�I�/%u"}�K�Έ9n*��_x�R)'G��b�|`���5r)z�A8��B­;|�z������/�R���*�E�~�s����YQ��1`z���]4�����҃FΩv��y5d����w�O���0]���^~�f W�N�G�S��b��)DC����ZL�� �w}�١�$����õ���B#o�*}���F�%a<.wQ�O�3PG�bo�6����p
 �q��	T�[��y��m{�|�P��Q�	���
�s2�~"�M[����ʚ�QA`/MX����D'�q�R<=Kҥ�����|��,f_�^ok)�=.�*�Էʎ�,5�̯k,A�F���3bZzTФ- u��Ŭ��K�]������>Bc\I{�JkE�K�A��"�m�lh��*~���BT�J��wby���F��R<��"�8�R���uC2��:��u_�Ć[H "��YT��?@$��.b�3��c��m����7��,��8��7R9�'�)��t<��a�cT�Ҥ��8�vR��wH�1;p!�����gI�7�H�n>�>�v��>}���ӌ�9����v4B��AFߑ~����l�u�	����eIi�굹(@�s�p��Al�L�'A���3������?���.�R��!�Þ��gG�`k�y2�O�Q���K\�I۸T�~]O�y;��	D!�x}����@2?��қm�2&�O�`�yƀVa�y��,2V}|�*�v�K&��6�����wE^�~�d��gG�y��SW��x/�s�&+�K�m{�0��ӡT�q���`�3�bZ�H������\!0	�`	ЂH p��*ܴ������H���n�e43�d�Di�y�׷pխX@]������d�_���~�mU7����۬�Bi�!���b��W�r_�O���ɯ��E�7���F`r&/ ��;����0Hm�͂mP��U�u1�9��!�6�G�#�6�ݴV�2��������<�E���K�w�*]a�R��'])��H��]ZD�+�{r��ݞ��h�\@Wa~T��	9ui۷
���a�_�(�+E ��J��.�����=��5ɛK�:���~.��	�� ��c�>�9�����ܚ�_Z�q���7w\~]c<�&�c3�7�VU�d��[Wߚ���i%��9k�հ���,s�>�ͥ�}��7�1c2ڔ|a
7!���ض���ҡ�^�$ �a)�z��4���F	׾��v#��j�z�����0�ޑJ���y�!�U�e����O���p"6>�bǈGĸ"7F��_�!q4����(ԋ�+ȸ$�)�*˴]�j`�uN�Y��H�@!���r(�pئ��c� ��^أ�����N��(�8MG���B��D��Q<�(�ds��]�S˂>��*�<�g�6��%X_�a�*�Y*��Y��{Y�᫢ �{w���ٽ��:���{�g�/8���P$��1 A~��������|��.vzHq�H/��*ʙ��*^�?V��Y̅&� �\����ʚT���ƙ_�;����N�X �k*/�s%X���ş*_��V����i�#`�����H�U���^u�_[v�i�֬�B�f�L�\p�TB�{��@�W����s��gmL6-��ѯ�3�4h~W'�lW�6�����Ь|.�h7���W=�5�钞�_�C�M��9y�{���y�\1����]��ܕ��Y�^LڞB�2��
�y8��p��Ո���^�����X��Z�6��]��:נ�n�"d�t��U��
��>�����"$jH������N=̐�� �!�yصQΞ�<0Sњ�>��i�mE�N�ls�س"{�	�G���}LkZC���<τ}kt�O��y�'0���Y50�1�g��,�Μ�'N�V�,��Ȓ�	tҸ ����o$��$��F뮬ݑ�$	��w݋z���ړ�eͻ�B�T?J<o����U��\멐���f* �@�����:G�� ���x�����ӷ
��@v%�0p�Z햌�+Ǭ�����yF��FFJ��Ѷ���TL=��{�ݺ���N7��Mƌ/��FT:fw4�K�h�xu�������K	�dkہ��MP�5�r�o���M��-����T�|�՝�����`4֑��f5��t��Մ@1�ɎS�*�Kˈ��Ij/�^���+\�\=K���9-��W��I�_V8���~d��= dmi!@�MuUD��`��}ҩ�0很��S��`���P��A���J�*a�xd�9k��:cv�# U��$�a���4v��a	K�G,S�t./�zO��!-��og}���h&�e�F�������9�Sn(l�]W f���ݭ�'�'K�\��9���@G�jw�C~^�+8ZZf�!��ښ $�0;�7G�$H^H�^�H�1æ��l����Ah�K�6�Ӛ�C�n��`�D�
1k�����#��Uz�,wu��is����dp,�8�Qbz��B�2<wu�y,���iʀ}Ri_6����F���E�����ǭ��#Jp&��ރ���/[ἡ	������χ2V��
GeK�r�	��ָ#�pN��&R�zu����w'.�N6��v��7hH�A�`~` ?mi���$���[�r��>��u>�h�rc��4��sFJ��rQ�˿)����&��n�c��>�Ҍa����F�ù�eĈey_.˺�V���5������Od`��m^F��cz%�p��ȸ��#��6 U_��f2�k��Bc���1�#��/�R4���������"a@g��U�!8&T�oTA�̏vq�Poc�\ޒ�n!����a�-C���s�Te*�q(V�K��M̹�wk_e���>�HkT4���)S���M�J�WQE�C�iyuς�4���8��^�[*-7�yTƱ�)8L��#,9sU�H�U�Kh�CIF��#����~pL=fg��kM����ت|��� �_�eT�c�*ՏzY�3�{i�G�VE9i��n�����CL��@!h[��,��tH)e�8���Z]C��s��3�c�z\}�l���9GQ"X싃 �&�#�6�h��An~��zX�6iѲ�4C��Bt'�	k�a��.<�ؐ���8�'gٶ�G�r����,O`2ڬ�1'6��	}g������#�b���+P�2N��D���q�yu��r*��sDk����/t�j2pP׵���9�iN(��t�E��� ��M�!Paߧ0VjQ�~�"�*r[(ߦܒ
̀��+�����8G���� ��G�1�X�`(��V�.`�{�X�,^���Ԑ��T�F�{ؽ�F�v��K9�@b�(���h�>p5f��@���.�XVb��̺���J�G����V�m�zw
L�м����?ӵe� ��ʽ����L�ʏ�q�-�v�� i�'�0����>4w�G�쵺tG����p��5��G��|r��O�%���ӆ�7���4��}zF��˪�A���y����'�jl�fu�؉�t0����i�����e$ܵ) ������X��Z�ѓ��/�z���P����Sڼ{���ϒf�y��| �0����O��A�3i�.�_,�b��ܚ������7�ɟ�d��4���Qc����:t	�&d��6� �XP���b����'��lNub9��[�t!��K�-�o��Y����Àa`��[�{�f�y6�����D�_��E�K=�3˫�q��!�F�;׷��q�l�(26�ub�>���tHJ��	4Ó��6S(z1�y�%�ojI�X��ѥ��Q#0f��,&AYx�?c�B���[	�W��% fWT�������w��`�	�M�r�so� �P9�����q�Nm��"��A�֚sd�ǉC0��	�{<����mW��m���	�B1gk� =b�z�]��^,�ԛq��%�'���LuNhJ�,�G2%�z|.g�$�	N��8��1@[5Y-*�J.Es�O?n�s���C�{��aE�c���bӖiP}���$Z"��:Ηk]���U��|�"���Ϗ�%�����`G|����{/J�D���a�X�3(Z7��DCG[C6j��
?��������!L����dO!@�u�f�wm]�k� 쎖|����18B Ň��G�mQ�*�^�'�כ�V�V){���湲�1�+�� �U�2�#��}mqӋ?��t>��ae�����������9QK��}|yN�8����J��dnN��<�t�EE�n����T�@�[�.�LI�V�=�$�аf�%62�u�P[�O���������rT���<�ߓ��p��+�`i�4����%fJ���{(�Z �H~,������Dw?�N����UO��������R��f�S�M�#�[891����K�#1#l���?�i�D��R��6Z���OB�Y#+�>7���ϊ���G�\>%�~K����"�},+j��YMF�d�!B7T$(k��Q2�%�o")ѪH3�0�F2����>R�{E� Vd�φNCԋ�4nj*ѫ0�I��NE^��4��Dh���_��Yn�y����/d͒���9���/_�4������i���6����0-��L��Y^� �UO�&��ϓd)��!|��um'�(�%GD��'{X�]�U��l��1�ޜ�}z�S�'K(��*e���m�ym��M�;;�jJ�~Q���YiQ�]��S��mn+���G���J�,�鴵��!�n2[A ��4�}���G�*�(A�T	��^�Է�ί�}���a�o��\�=nh�7
�i�q|�����K��Q����^��Z=UFD 6����iQ�����Z֘
 �"�>\	2oh��yU�懓*>�q8G�C�����Oؽ�D.�e�RfN�{�C�;J�j�#�xv�q��R���� �3KP����Wh��K��a�-)+d)�l�\!�6Ni��R�E��
K6��>��\�}O�B�Ogv����w���F�h*�v�Sal��J�[G�u�^�晣�������]O�.�M�7�
���%�0��ڈd며����K��V�����`p��5p<�Mxv^L�o������sdPDn����uA9��]�A��w��?:��S�]�M���_
���[ʱX�����V(RdR��p�,�\[�IaV�9/��9�lқ펒�nCW�d?A���`v�L�4����J��/���  �����T��Pիm���|����2�{�$���4��j:$��.��ß�f����M������cvfXQז�W��(Mou�J�
-s�����JЎ������Uu�.��q�0F�����A ��1���Z� 0�PT%S�ڞ<�Sj�э��2�P�ăoqǋ�yX(P-ӣi�KT�]�;�=�456N�(Aһ����\!���w��$>i�z(PH5W�jh�;M�BolR�ӑo0�J$F!u~`K�P޳��]����!8�ч�Hsu��6�˜��z����Q���v#��N�';�*[`�o5�n��<m����?����?��J�0�θ����qcOB,��6U
�K�5�y�^z���I�zL���mٳ�芠P� V=�@hf���#~�:]���s4Y��2��ix�Em1h�q~'ɔ1�3X�o��	O����*��
�[ �x#A2��d6�6���y��%�>UBs 0�S�nܑ�Z�&�°R0Kߏȃƨ��j�%[������L����z�嶚3Ӄ	Vf�<�����������j:à}���!���)�g�8H�'K�u^��8�Z&��`��gKZ� ��%3⹝��|�p۰}31M��Q��|�Zj_H�gS����I��GA��cǈ�������sQ�B�x��ǹ�4k�}y7T���OA:���sҠJ�<u�l�K�����8dH�����*lM����S��4�$AuR޸�Aov ��V���X\�Ꝧ�q�X��3j�n�
j�o�l,����B���ա-}L� o��P��y�B�X�`I��ܴ�^H��X�΁0��M����SbnL�jC!���dL ����"$D��̀����O�͈IV
u{a������{���k�'���d�I!����n������">J1�`x3"�Mf�Y�7�D�0��,�� AL�g�c�(t��S?�?������+W��s����@
�*�$3g-��B��5��?����A�~k�uj/��7J���Z��?-*p���s��u��Eq�����߈�%�ڥ�2��~㗀S��^eo�ި4
F�{dE(�2��c.���4�;��us^�z"��4LD-S�阑xw���x�:|���$k�}Ԩ�V��v)[H�x�G��DB��~3f�G�����-�J%�V'7�x$w��/�q?�$��)��bߧ��ʠ/���-�?�WJ�1�a�mJ�@���a�rP�&�EjT�9HW�K�T�q��7�����r�_�6�W/c6E��a��.#p�p�*:���t_��^�*P�NfO$!7�;U_`����N΍�٭C~ϲ3Uu5'Sz�q֓��ⓜ��F�� ���q������JG�C:U� \�����dߵ��W���!����r�G��V�o�&���2���9M��]M ��1c[�¹�H���0�y[�=`8l,�UQq�`Yí}:WJ���,���O�&��ֿSA��9�OQQ �PJd�R�5��E���>�w���.�3��o�M+|�W�\�)����
]E��/�,�[&��n�A5�&��ĆB,C�SX}Զ�~LJ*M��C�l��̓���A��ȅ�"��L9�����j.H���Jn�G��^�zx0L�Nw��n7��,ܵۢp�9)đٜ�*z+�����p'�\gr:�����}i����rn#�BT�>N�)O~�D]k��#�p�ʞ�^6��[�����fw�➀�z���y�+G�fӋ���{d=��N��t}�o�I��v����s�r!�cM���m�5Ht#1���T�d����ۣ�!�{�j7�7\E/v�|�/�\dL����Z,����N/�0ͦi�Pf�k��$�ׄɥ��b�N$n�ܷ:�7��`�I�	���hD��V�fg���$����Z�%N��'����^��GSly���c���?"����y����^2��~��g�p;��x�4��>ݕ��b����glY�ЭD?���9h���X�
rj`�T":�����P�>����{cH�/6jA���F{�=�%��[0Ȟ���N��Y�G%@���Jo�Zs?�B�/�2�W��PӀ�Q��wRz�_2mn�D	P{� �,�Zl�w�/�M��X�	�T4)��t�@�6R�H����������|���k,�fxl
V���)�f_M��&!�ޓVl+�2m� ��>B��-YEOM�<���P�F2ڿ�����j�����Mh@9`c�Ip�M�sC+�����0 Sp���S���R���c�We��n���(��d�;��rSo'mR"�b(C����1�vXU�I��I��@�v�����p�K�*'�R��88�%�N��^,P�=i������*��\�JiH<B����C��m��9��k���&�s@��fB�?j6�����9'��|��Լ��ٟ�5rD}d�x�E�;K8o6�ۏ���K�7�+�A�2���6�[V�Z��l��T|� ��۸tO:�K��B��6ÎL=�q<p$倬���?�w�JIo����}�xS������c���W���c	��4�����~4��QS��ծi��9��>��SL����)��a=�!�2�e^�0=8n>�2r�#��'�np�A��Z����?
n6y��E�� �a���G`���L��F?�5U� �.��B
�*F�3�����Cy�x���L�x�"�Ѥ]��=H��w.�`��z7*��`�K��<-z�;��4�a�+� ��䊻����Q8���t%`m��"V�@�vc�j�|��y7	�R�)���o��ؙ��`��C#�>�-��Y��4n���"�e8ٍ��ks���	�x�����Z��ǉ��![pɶ�D���K'��:i�<��2���)�?�Od��-�G!k�v��n		\�Z��!?��	I�*x'��=R��D�8����\g]����h˻I�G�{f���[�S�u�ĩ\�tY��Gwc�@�"\�M��J�Aw��yℹ�d�]5����<�1s F��;�7-ƅV�+���N�ش�b����͔����摸_PLWƯ����.��C�L��04~�$ۃ�(��/S�9��!�����I�N�N|B'w+18�_kx*��'�a^�{I��o��.�B@(�b�u)��ʢ]:Iq��F:	�H��������Z��Vƪ���'�=H�_��.��w�4�c�%rS����^k=�Y�ۣ��Ҽ[�=�;�j}����${�I&9��֫���uJ^m/�(Y����^�8���N�Jq�"�e����(�-��߬�<��S���y�d�H!|�)�ǳ�m��ڊ�I��RBF�S/�9K�e�?/�=�}�~f%���{m�#�	�q8h�5�D
bz�[Mo@Q�y�D�}'�*�(MV�E�᥆�g�S~��T��P�s�j�7�S���b�����VX�Eݔ�����w�,8qU5��Yq��׷��0DP\��r{���~e�%�j/�rp�zP�W�魨��ͪ�
;g$Yf�U��g�0B6�;(^u��-l��� ��#�܎^�����9`�\�0T�_��>�P�ݿ"i[Ҙ�7����r~�Ѣ��?��OG�ɢA�Cb8>��-�,'?�}�Q*��.?;�t�>�-ױ����>��-�@'�7��7R�&2M��ObT7e)6\�O6�pO	^����K�Y�Eo�Iu�D�:�T1y�#:�x���X#�YL���U$i��^4z#M/n�Q��Ч�"Vqp�2��lm��A�j9@�$*�<�b����_Je>mu*)���5�5+/[��Bd�E����Vx�M!
�F'�J�Y�è�&r���8�lN�qąWc�Y�v��2����ЩrMZ�S�q�����G�16��&��k�> �0��dP������n�����!
�|z� &�(�q��_$�C���"�̱V�H�^R�e�&�9���ܠ���z�i��ߢ�x��.�v�F)��e�]��2�D�_�h�,�����'��&(b}H�Cߺ�Uk>�$��
�7�q�^�͡������5(������kT��H���v���b錋��C��l#�9���TB��S�z����`z~�Y)G���AH���2':ɻ�Æ��b�Dx����#�ِ��\H���M�~���CSI'��4pnH��,GӺթ�D<ԘG���R9@����j��5��}��=��6��;�!�yf��Vt�������L���"�����8ѥ�j�7]��u<4�r��#�'��Mwr� y)�+���x����¦���a�,5B���u��~͍:�j:��/�� Yn�j�����%��:Y׵h��I<هx��Sq��/��4B�'�3��".�
��Ǧ���#�=��'���@x<���@�wz�����T�P5!������|��@���M|�ԝ�/�քט�.�?Ga�iH�8m ��P�B�®#ݕ����3��Apb�@�Q@>_eQ#V�����q'jZaU��A?�����zϟ�Q��|$��,BԿCJI��ך�@Pv��2����-#�PC���0��Z%���E��B�����r>�	@�I�m.�l����}�(d����O�i5�G��FR�osU��#\��=��~1�G	�&�Ӳw��4p[�4J��J�S(�a ���o����{��ꂃ�%��Z}|j<O$L�� "!(��rL��Q�R&EuvB��o�'�� ��oN��T1�"T<:V���_N���JLd�C&2řY�6�[�p!��@M���@).����ٷ�o,���d{B>!�\��Z��5gI0��U_V��A\̻��k��N>y��Wgm<5�T\�@&,�܌���)��~8�ćn�H�`� H�@���r�O�XK����z��y���̸�:qR���o��G�Qy/�i�z@7*�3�\ҁF���ǔKy�����ttk���Ye��=�m.ֶ�j"�}/esj=�lU}���F:vR��P�T�4�/�>����Ԁ҂`:���c�H��+"�`�,��AL�Iʏ����D��BpLeT����)��JQ�qu �̨�>Pypl+}��m^l��z�;�e��! ��y��k�!�T��~��NE�g�DA厈lR���3�{7�M�G�Ik<��#�~q�TToE�Y8�l�_t$��Q����B� ��ub�1��t�a���~r[�4��}�[��ೡ8��O���n'���\z��D�E�Y���ۿ�z�x/��(xU���B��r�R�a�� ���c���$�L�z?�揲����Ը�P�~p;ax+��T�1��S��
r�f_{��C��!M���zUD�$��6C*��T��H�W���-��IY�uޓ
�����Ye��Ti��nZ��Tx�����޴��L���@��QRn� 6|ŭ�7M��GIixJ������dWe欼<:]���N(i�;0�n�D�
w�4���l��c-T�G���xR}�ZC	�1�%�L�*Uϱޟ�7J���8(�~�+�Rg$Z|k��%���t�H�n$�U�ʿH�S�����H1�b�>w6�K�P��� '�AWXY�X�8!]��+Z�|��?�lD!N�Q� /��A4��X���G�5�,���g�H�>�a��nU�
�W��������V���M�b�&~%2���q)JA�#��"Ie��C�5��@~%�.j]���?:��~ƽR��F}  ���E)����^B�~$���ˌ]N!��=��s��Z'b�L����Q�YlwLl��S��C�#�m B<�� �P=$�܉O�k�+�9\�.���_&ИH�!����RGcuM���{����Y�o�������=�F��m	y���J����ʈ#\�7�.a�'g��"�[!�*����$�+D�ۅ�k̃N�2c|� �b]�[�r���;�|q�:{��774<w)��T7y��%c&�Xc\å���fI��G$S�1&N�������Q�f�H�۴5-��T��n�|
=��'��n=�O�q�¢�Wn7�={�&��!W���hv�}�<�4��$��;��,�[�^{�P\����s`�Ow�i�c-o�AB-����bQ5z�fY~*���i��@.���V��_Flz����~�bُ�D��D�ԭ���������H�ɞ�YO���x��T)=����I�>�8�Y���pSgY}�'�h���R��?�	���v���*yQuÄO2ف����̽�����ױ��c�40e:@�Ԉ��;��$��܀�h�4⛃��i�{[�Iݑ��%�É��7�8�������V�k$���j,�1<�"�J����Iڽ��@D}aL�ki`z� pߺ����0�$
Ax�Jy�(>E�����.�<�G�?�A�%�͑��?��W�D���.���;]�x�^"{Asw�gC����2!�F�ľ<X��5褺9���3�3�SK#5ً�%Y���0�CM�x���-	��;r?�' r+�����1�TE���S�����]�΢~�%@�<"j�=:��,Ч��?���]���uR&q�s-NAe�xYH:N.* �����1y�2�<6�gѕj�#R��� ����&�m�h�	T)�V�a%s���U�?�3�	�u�s�$ҥ{�o�&�G\r��	�ױ��ѷ;�E�]��4��C�1�(�������UF:+�i��p�C� _�oFUڧl��W 'M�g�<X8�'#�;ۮ�!�^��<Ș�I}���SSҔ[iK�K��,B���A˅,S;��)nՍ��>���W��.0�l.�1<1������5��s�����5�[T���|��$��ݢ<��^���C<�Q���vM�H�]�Ճ�J5���4�w�Jj���s��H*ӽ� q| �^����0����N�Gy�o��eo���@�+dAz���~�3RZ�������򟫲��4F��S@j{ܘ�[�$E�ɐb_��!��`=����Y�����f#MRS3�/v�MOJ�{��N��8%B/����VQ����
�}b@��7��(�����_�� +�M�X��/s��V}����B��4x��
B	)���G�oI��媾��D���q!�3���4Ə9�ݸ������{�E�ɷ�6��g�a���.�g�EA�m��"�zf1]�P�N>i�<��qD_t���n��mV1�HF���x��4d�џ��& -�n�Ӏ��r�;'�,F��\�nސ@�vG�w��:���+�
at�X�]�]��������c:���wJ:�խ-_����k� ��J�Yo_���� E$M�$$g���*�����y��f�����	z�7��9=��r�`D<#��.�1f�1�!y5m*K$�o���@L�S�8ΐ�_VFK���bwʤr�b��="��^+8��'$�s�9Kc����u��Qk�>LMs����X�Jfᔰ�l��F�M�HQ�͆Xl�^#�N�'C��T'�^t��l�Z暪���v��$�Ĕ|�����l��+�*?�ltL���'����o^�ta���C��@Oơ�A���^H�2&����b���d��bi7�����^{�G\�c3Y�\Il�F�)��dO���b����@F�oum��4��F���_��x��v���=cIƲ6��ڞ�fr�ߍ�Dв�Ł0�M���C�?�0B�_TY��F�
s_�����;^3�g���>�-[��l[a�R8�>�7�$�3��{�]��-���=�c��%e-aU���/��
�`=Hfqfl�ʉ��������B��*�`#�$�]��ƶ�n�!�U%��t��l޾���絆�eS�����%E�^�xjБ���H�I�[t�`3�z�vX�gsWg%N���fh;?���B�=��Asx:E��oQ1��טb�O�F�U,d��|$�S�*�.:Ã]�&��Coqϔ�&�a���*`����ao�X9�M#<��~�s�Ƭa����~�fnmQ���;�h85L��^"ݡfǧ�gg�/��U��� S�b�%{����l��P����r�l��L�ʚ"Ѝx�\A|ڮ=���)&=km�����w��_ D�{�٠�nH6ā�=�Đ!��'l���[Z�
��$^���mc<��bX�&iw��J�EZ[��>�^u�H��}�@c�����$��(2��q�Lv�RAz#�'2ӫ#=k���`)�q���X��1i�U�{fc�����ځ�6�JL�B��##�̸O��Z�����YK���w�靉Gv�g;��n->%i��ChNB��@~��k�=j��S 1ɕ�kP�8�''Dޟ��vmJ�0�:6�*��=m�i���&q�;h�=�ܽ=��ox�x�c��2�n�ҋ;�J��1^:�BC>�K�0�L�1U��J'�߼7�g�}[��r;�ࠔa������#v�,a��	�O-���6��9�*�ТNz���E�/m �u��R JB=�R7�@��X�T~A�-���{�S��2�ݫm?~�k�؀��tI�ۜE���y�TV�D)f�dskX˱+��m&�\����5���D@�U��n^����nn�\>`ٵI1�-�w�2�Sbѫ�D�b��Ḥ�3?�_����F���RW�\����j4����ŀӣ
�u$|���wJgҾ&�)�?�N��n�{�%1+���������%i!��<�}xF��6���L�_�a��Yt�tj|��JQ���^�����ν��bo�M{;Ն�9ԇ����^���P��lAL���i����j��x���~�|��챐���gͨ�_��h�O�X���t�S��ǥ�{s���8��-��v@�\�=C`'IJ��c�6���n|1�t`MPc���m����~�Y��%��J��=���� �\N�������l�y�}*���(}2�|6HR� ���׆wgV�ml5͵Y#l~�l��lf�҅+�+P��(�0b���ǄG���"�r��nF�B�ǈ�^��L!��GB�=�#�q��FW�[�׊>� .�'M�Rx�5���1? �s9������L�2Z}	e%��l��'��\�U����jP�٫���ۧw�Z���=%wU��1�,��>�dj����vBp�f=��4׹�����x�id��Lu>�H'��T'7#Z������^.[��/{�	� ����F��_*���2]i��e@������]��Du�D5���Yd��%:ɼA6JT_4C�l5v'm��vU)�X%Z����-�l��2�J��[�"7��?v�/{l��}�}��⿲B�A�{�Pۛx2��V�s��g�?��f1��- pQnp�V����_��������g8��b^��6�K� 
N7�BX���Gpb�������v^&n���Y%���}������S;�m�H<��(�M�`�}�1 ��A��[g��	�e�W\�������a�P.�%��͕҇ T� �au���G1&[��C���|_S������S�*��������ַ2����+�L��R[L'��~�r(��g��l��= Yg�ҵ!�3�}6\Mx�e J�c�x{	J�s��8�i�At�����~P��8n��/z+��V�	[���T��v��5J]^���=��rzG�?�������2"U�;�#{n�7�%r��Hڒ�WL��=��zf$+줸du�<R�P��-r1��e7Y���	-�Tc��B�Q�"A��e!7��o@�#3W�ѳ3�˴-n��?�0��2�j���
�~95N���@n�Q���	sGaW��i7���h�Qf��8eF��m���FH2G$�+�zx�oTd��I�l�@�3=�sVp0��nY�����<v%d��oq�^;��hx�0�7�9�e����A�?Y��R�*\�d9�(a�.3�/!r��w�����L̊�^�%��,&�ו�0)z)�.h�����K�5�)vS���!��Oi��sx>���C7r�N� �C�L�8�T?d�9T�dl�;�� k�h�M~�;g���2��G�ۣEn���}�lp*%��ChFu�t�f<��y����~�v#�,�r��-ks���C�A~��EB����r�UH�8\��p�I�Jq�S�C���1�0<U3�@ ñO�Kf��2���5S�_`ܪ��\	�Q��fl&�ơS���<�Q��(�a���mE�mH��z��W-��sk]@W"�ߐ���(ԃ����uP
zB[��4^���#���NNI�[�}��F��|W����W0ِ���pv�I���ސf������B2�{�.y���(�C���j�YC�0I�/0��v��,ܰ�zEd�+���Z����$��� ʉ�,����)�^�
Ң;3Q�q�(�OEl!*/P�iF-�����r���,<�F�i��d��FR�1l��j������&�����nѿK�W�}K����G�����9������=������E����hJ���CnP���?Q����J�-�!���+!���6�q�+���ϋǜ�V�/j�8���57ƶ?q�0��q��	@l��~����+A��נ*�t=����_ų��إ��L#���!�ʂ:B�?sy��ת�Շ�2{I��cC��W�t��E���KZ��l!Ql",��X}�Ͼ����_f]yh��.ဝ��L;@��Sq���2ҼU1�M��g��DQFMgQ?:0{��4�^�P��#���%�D��&����;��,-Ԭ��x�Y��x��q�2Z�-��(O�W�۔�$K�﷋T($��@��7~F�?�֝�ɽ��hP�=����_Ygi}�����,#k��2���U������}S(S��#�u����~�P"�1�\�Bf�=��N-!ZB*���ٸt໳�&��z��X W�(�h)�	W�x�Ӏ�����涫gNqLY�;�prl7�q{S]��s%M�7����g0����l��ZЮ�%��M�u�K�;g�,��@�a��
�n8�.j��1����d߳>�0?$z�A�S��o��v)-	4�oJ	��{���n`�R��ATj���i�����*�Fe�ȁ�Y��{5|�<H@z1v��f7�R��/���&�
�3��@:�\�6�9�t���7&��<s��,�4�Yy��y%ܴb���G�Q����t�̔�k.��/�qE,�A�����U�l��cؖu���'��	���ʏ�-~+�]Ȇ�6h��W�ϗ#7���[PI�[〈��<�T#�2b쯟e;�kF_���s83�FH@.��{� _�Z�j�<�&4�g��<�1��5����ǐ�a���n�G�э&#��h,��_y��t޼9��������=B�sO5ѿ����υ�#9�9�0����3�9~jw�p�;���k�$oQ��h;�vɀ��r�v��:Z����|����P{�FV$�Gʕ���l�| �b���7� ܗ<���U��<�ԟ����\�`4�mT ��N{}%��{N�I*V���g0{$�Π%��?�;�3c����k��k�v�)�4/=�f��A�]��t���U�|j򗺃�T��xE�sD���c�?Ǩ�#�?��O�׾oI��V;��iP�1�[T�rr�:���L��J�m���>�k�1���| �ں�'62�l��j��Gf��HK�\���)���H�7xl�T�UPi��>4e`�d�`W�rg�2%%k��:n���g/b~�X�K��l7\]x<9�z�..�w{!\�,N49U�D�?��W_�q�M#�;��ā�Ig�{68�b7��y=��	���&��>�x��981�X�!��n4ڠ�;X��Gt����h�t�{m��GA\8^��ޥ-M�?��r�#)L�7����ב� �W��\�܄�)eK��� 9�&��G�F���A^˳�:�B�,AK��(�gЬ1n���|�Gݪ�&���}"��u�g�J�8�B�ՙ�ז�"rWY��N��'�0�_R�6�}f�V���2w����N�M!e�����D YBj��T����n�vV�||�X��p��5|��R��G�s.�qe��R�
h�">��˒d���9������L�>Y��-'R0��v���"�)r����h��N�6J�.Kc�A�k!���?����ĺ� r�Ѭ���.��0U�a�Pb �`ZPTm��[p0��r�-�|#���fʵ�D�)��Z��T ��&���_�?�,�ݢ���5mx����j����W��S��S\	�3u�34?p5���{�j��e�����[�C�~[w嬣���
�H����u�ȕV�?�$�[-&b�}�Ut��_Mn�k�I�h�=πF�᫻tS���kA�鍯;���]?�,/RA��~NWJo`�!z�.l`��)�����
��C'�J�����e��OP7���l��]�L��.�9l��~�ǡ��=�֯Z����V���B5>�}ߠ��֜p.r�j�����\�}- ��e]��]t�EF�|>�m��"�J��=%�/4_����W�<l+R�P�_W2�j������*�=��ZY5�#�Nq%�Y)��X(�B� ��Z� ����Ō�P������k��z�:=�D�2]��N:�~Bo���y�a��UAOʍ~��=�e����vW�+��30�-Qwil\)}�pE���'���{�&?ft�)ߦ�h�g�g>YB?��-�(�*�IӢA��.*��#&�`d��wA�;N�4%.�&"���S�k!?��=\'��*X(H�j��0�^S�&���&9�_��@��TnQ;��nr)� ���P��}��\�go��nk�G���Mj_L���_b�v���H�Nm�֕���H��P��_����'j���<_�^U	��M�>4�G�;��üh？V�{��̆��*�2º����.�AM��p�hg��%�T?g�he�ٖ��k�WD3Y�tL:t�Mvs�)�C���	�W)�+k3Th4���|� ^|�E%Y4`�������,�\�l�u��)۷AͣR���'0X�ӥS�[o<�+-�(=*��z'��V���N؅�S�P����}�`9�ʟ��O;�1mAOnv+����D�5(:��	qg%�ርjS����.��$���8��o"�7����[�q�VD�ƓF����<Ip�h��?��x)�������ځ�I0~��͇�ޝ��33�oy�<^Q�q&����׏eЭ"�Ny�d�9�T��+ � ����:��ST�!h2�&a�ޝߌh
N>�^*���C�/��0J�\�t7���Q���R�&�r*M=2%6�K�q#�l�\VH���ߠ8��լ��Es�G�OՌ�x���
�n��$�HW�|$#9�z�@ �Y�/w���<0���?�b�H'#��4<��H�f�e	���F�U�u��M�r1��,갚���I-�Z�l$�|Z��Xid���;ۗK�5�@J��������AA��oA��s���p��cӧ�ԟ	��Z�r�dhjB�8�8�����e�E��r�#uO��${g��RkR��/:��TVq@p��7�[z�γys{{ZH��Wɝj��0�"�y�����'G���⁝CakYl�i�}�z��Nد�G2��i �~�Ӓ��F�D�'�����ɚ=�Z�t���g�Z\�˹4<^���;�c�,�޽˥(�@f	��i.b}�ذe�cS�:�
Z/>I,�������(����\�Ů���%�e��B�B��0�G�� ��#���/�?�ƈA���w�W=�f����ɤ�Z�gߌh��y J;'G峕T�����&7����"��M��,�}���=g[�#����P��)c���^�#[�qCj#���y���T`^�L����q�qQn���<S�{�>�_��܀-W�f�lUeV/)�atD���f��e"�G)�`1�#;�=�������y���/���H�d}()ʷ��-�@ ��yT�p�J�G��o��_i�K����S7�p��ǽ/���N��0դ0HT���"����aA������"��a,Mb��Ȋb�@t�nU����a��W(�C�<�3�R�z��Dz���\hR!zc�:�P��X._�s�Ñ��y��ؘ�7b��
�0wǗ�	�am���9T"�(u�&|��ۮR)�J����^���G�a�ܨ���vk���A�g7�	a������\j�S����UK�WW<$#��f/S0� c����r�V˞}�$�(��Z1Ӽ���*��wg¬��P��W�KY��~ጪ��VY�7K2�JjM?�x��W���=Ρ�޳���@���[=<���j�}��]�Du`VmV@`^�&3�i���^[�$�-��}k4[6(��������ВFM?�1b�g�Q���L�Mi^�������8Q{AT��h;��6[s�����7��ţv	���]�
�M��q<��\��5�W�m�0{.�S0��PI�$�!`@'�,@|�U�#`~�AV�������|�7�`}�@ҝ�h�h��]C��kc!������~�̕����eIZ�8���ɑ���m�A@(s�.�@H,p�T�NA��fT��6����1X���h($�s�7cJfiAЏ$>�~#����|�xt-�C�M�>2�N�{�LU�c^nI,clD�a)&n���\QSЎC��Mݰu|��;�����%��(�FT�������[��\@�h@$�^K�&������Đ�ۑ�>A��((׆���^w�p�H��Ϻ��-���`�h8�E�.c�UAG_e�=�9�C�K�9o��b�cF��P�]�_�*A�8XPp�վ2�ޯ�5�Q���F�$v�^��{����@h>���k�kg����&*Zh;c�S�Y���KA�p��[�1�9_�`���N�hH��tsoJ�c|�J�������>1o����CJZ�3F,<eƠݠ;�a�W���q���L�f�;`E�v��$�/�fe�������S<.���ܲ���S���C�rD�>�̾fX��oVjaB��ֹ!�)��=1F���e+�vd9�Ig4(S��jR�(���%���3+��P�7�yւb�6��G�#�QѳfZ���"tD1[�Hv,�9�(D8�*w�?���)�d�LR�ȕ#,��ڻX����d��;����Y��MgkΖ��}L�0��ȉ���W^@��!|;�M���?�)���#�3Īo�������,Y�Is���H����2� $��VҬ<"�ֹd"�z�0�ٞttG��}��B����@�-�����_I��}Uќղ{��-S�m��W�qRS{Z�{x>�,�:T�����.�Ha���o��.�w��R���<�̷U[��RRD�p��Z�:2�I�V�y6^�e�*:��MlsJu<$���ٴ�;k�:*�̕ iy>���f��[���[V��.�:�u��sR'�'8��^E�93
=@�^��pH�_F�w��������*�66�����@5��(2����לM���P�t���X��������t�������+���J�#� �rBE�*oOP��bp(� 0���'����
��h �M��1z�Z\ƿ��]���|���l�X�4n!Xqɰyd�жk2��.[^`l�dI��JN�_�-hSsۂj��"������&*���	���~,@�O��i�6)	'��]w��X�ܒ'}��%��F���P�>Mm�f�X1��ڃ��T#��Jkt����W3�U/o)��R�[����	ɥE�I���7d�adÈ�k���T��B�p9���@q;ͺ��} ��P���<��k��-| &���A,��?�98z/�/�@�R��B� 9�C��� �ƓC�n�%�,���h�Uw$�0�7�P��2�Hqó7�ՂPL��1��eq�<_����0e�b�2��C������O�Xk�S�:߫���R ܞ=�D�?�F�o\Ϟ��⡙��o&�o�&�����p�:{J0?�R��ts� �:�^���s���NL�8�u�f�A�MN����jb�ۄY4_����&���u��*\8��ksH��-���1�7a����mX����l;!F��~�p"�9GE��fW
�o"�'��ir_�;w-�Ĳ�� ��d}��"�;�C��vM���9q%t|�*�-�i�~���|����bE�*���M�k��|�b���Q���l�$a* �2Ӈ��yz!�C�GZi����c!w�1����$w�c���
����P�:���O}_�1�cQ~���g��"������-�Dɖ�^�"
���1�
�m�?�P��u�4�=mq���[�[�S�!������)�U;��;ư��E��V�t�D���G�'բ��ٵ��H��Eϭ�#���(����lv��J��g�#+9�!!�,�����m��IȘ�us��d��J���oBǌ�u�T(�vy�p^�uC�r�%`b�o��s�O���pX�����L�r��n9m��I��T�����\������'�$��BPg� �1�U�Y��|ɋH3���y#7����Z��,P��:o���q��v�3�M>����mޑ	*6�������M6���ޘ��)���� 4���ʨ�o�%�[��J� ������9 ձ瑲��}S����頋�@�$����b���T��Ƹ0��5�sH��V����I]�J�Ƞr<��2x5�#�P����;86wO)��~�	���@&m�eAfRӻĻ��PV^��
+�H�Q����i6���,���T�L�r8(�z���+����#��r{���s���WbD�lϪ
��K�O�:��GS�9����0�g81Z�c�Q��1ä2�"MTN�}�-��0��rJ���6 m�#w1�!�t�UGZ��3�J}��������ɢ��u���mJ�%�0p�*���P?8hq �y��U�$�l�T}��� x�����Sl��Q�1�(�?U��cG �����gZ�#/����|�����9n�9�۫3>��<�����JC�<��Y�B~���� 0��;̗�>�d]��Ёh
��EX�cnI����[d��BЧ��@m��g&h06z�yP���!%�ꢋ���}2����{��h���G�ĩ��h�],ڃߤe]�^f�'�=`0�ʛzb�F�6W��.����JG���;�H���s�0��������%)6��C��Q~�j����( ���؉^��׻/N��
Y�ʣ��j6���@.�Y�%3͢�ϝ��4
��R��/��N!�n�y��Y�%5��-E�Ѡ�lD��A�#[5!�Up�����)�c�ƽ/��qӹ��gYjJ�!uʧ_N���!0s��Y��E�\�`�S�uu�bF�8����G���s
)���[�E�9z��i��
�F��K��f�]p�������&c�6#5�H����։�ogX
2a���o��!i�[f��o�(�� CP��B��b�\��k�ƺ�E�EDe�7�N����h,EV5kmyi?���np����yڿ�jƪ�o:q��䴰�"J�UQ��\�T��
�#���y�n�µeس-�pk�Nc�$v���F>X�M89�B�E���\9/궴��P���`�k;LQf��F����b�Buqv,�c�.N�#���Z��9�\����T�l��rD�3T�'F7�-�^Cv��p�D��ۨ~����7�(7��AP��c__)��u��z��%Q�GG��J����>{��k��%E�'){LQl�U�w�|���9@��{U�%�������3��-�/��g}��ڈJ��0HQBz�ŕIs�:ټ��`j�����3�������,�B^��A��[6��{����"�B��hV`�֊�`��vU��]�� Gm�`�a�CB$��s�ײ�V�%`b���Ў�+r�J�l��L)��j��4�$Z�0�k7�����*�@n*����aa#��t�y�9K��V��yBه2gݧ����	��#y��'�BG ��B�-}V�|��c����{<^4X���9�M��JL��`9�<k[g�?�����B�C����ۺ߸c蹷'%���i�`�K�W�l�S���������l"q����m�	�\�g��Y>"��k�����\�
�xH�=iu��͟y���K���3�y��YS��h�.��Od�Jj�T�Tkm�i������8����w���Xs{@/��wFY�x�{S5�lc�
���4�Œa��j��#����Sc��C��je����?�Z�-�jKo��H��Ǝ�d�^����w��-�WV���4���h�B����]����4pAME����396�H{�V-2'�u�� �� "�fb��:N������Wpl��Gc$,"�9VU�q�
��1K���-I�9W.�?Kɳ���6��*x��0��mߓ�,�0�]�:`B馗tt>�'��: �-����)3ϟ�w�Tڎ�m`���Xi�~\���{f%+�z��?8>�Y2������w�c����f|"NƠ~VWS����Qte=h:b]�g�t@�?(D�Pe#��^X;��P3�v��&�-�X�R���u�+�{ܲgC�`o��b����/v������{f:g�I1=�\r�O%>  j���Y�25���/ۨ��2��}%������m�"�k0�^ܸՄ�e�7���^B٫���p�@� #.kW���"�ЎU���dM��v�����+��S�a�CU/�/��qn��vyb[�k�@�3y���
>A��G��ӏz[�R���T�i�~҉� }̈)�p�6q9�A SWT�u�R��$
����Bݫ%;�j�w�2gGi��M�S��Z������EBq���?��|�a�*(I;������^iHvX�;�ld���NRP1؅C��Q����0d��`b�NVx�����}���d�ui�9�H�uN���T���#��ƿ�ꀬ�
��z+�'��0��6��9
T ���~H�2׼��쒌6��Iͺ81����EI%p��.�'ch�d,h�U~ӡ�]Y��,�w�n��=��7�{��a�UBc�;�.�P��a�}����,du��M��-`����j{Z'�`a�1'�II�i�egc����J1�C�@:�튟�']
��t|�;�Aa3qѧ�I2��Mz��+סYA����I9~��Ԗ{S]�-%�I��p�B��� �)���J��Г���V��m�n��t�y��c���͑ں�ZDg�'.G�h/�ؘe�ʁ|K�i����6]Q
�j���d*�w�8���#�C߼B�lv����-�-�d�<�.U���y�Z*~؂qd	�/�Ҵ�3r��?�K���}�,�*0v�x���"ȩ�=�Ыb����u2�"�²yy�Q#o9�\k�,Yc�k�U���;p�㡿e�uW��ح7c\���),��m��D^PƖ\�&�%�
���)�i��f�����L�M���ʫk�)��W�y�NmwO/�����F�m�/#�/d��i�n���I��Yu��fJ��T�~.��(u6�E�f���f�͵�[4���W�,t2�R��_.�&��<�b�G����lQ�9o7k�vϲ��'J�%�^��}!aQF��\��sd
	y��^z��������^�Ӹf�ʉ�DM�[b��x�,?�DBRI���1@=c�̻s��Gڂ������FW0o�pJi��q{!6�Y#i޵5��!Z�ݰ]w�n����`��ƍb��,L�$� $��������|F�v̏����>!¶�y�����D�������囬(�ӷPQ�\���|�"�W��|�b@��C*܈2ۇS�I���X�!�Z6q|xc}3�v�u����s�B�f���T���ӹ��
}K}`�\�Ź�M�!3{��۬'�Gi��W�Ff�5�_�f��'Ȇ�ςk�6�X��)c�ĕ�`�.x���.'l���V��|����M�矻h�R��ދ���=��R貥��#:�H�E (��϶���#c���h>0�ȁ湍��0��j�H�u�/I���tf5�`�o��6Ĵ�-�ۆPm�m{l�R�,�R��} ��:}��ft�1x�K~OϬ ���#��hk5�v�X�AɢG��=�>}�;��f���[7oU��:���xm4�����3~w�O���?t��&|�`K�a�slf[�ҞH���`��@����c�9,_�#
@4(u�K>}'c�T���ɰ�˅}5	�U�S��1`2�J�V��|�"nL�\w� i
\�����ײ�YQ@Uv:ùG��+�*�~̤v�y�.�;�'��:�2�-���q(IQ�����צ6�j+Q����#3���Q4�34� �!RvI�J4���X����,ƿ���"7�Jo�_N�.�@S��Ȉ���5�C�\��v�X���G�	:|-��|"!*�c��*�V��8U��aM�Vj*v�*­�b�n��5tװ�s�݌n�g ���-�~H�i5��c�%�$~).Fd[@A����#�rRH\�����|�*��*\�#�E�1��U��.�4٨�ψg ���Lf�hE�+��$:Bq�%����\O��gw��2$>�N��W�U��A`���X��Q`�b��h�����ggq����ج��|��4s֥��!����c��K��R+��5�D��`��Kż�� ��S�?=O�A]Í^�'���]��H��-b���� @��9���n�N�*#�P�����\�N�h�� M��k�h[H}B��$8��	�IGd�-���B���~�%�N���b��HI.�����y�;a�%�ڍe.e)��"^ۧ�:���:�(�5�d��l{��=�$@��f���K�U�*����e����q�S���e>�ظ��~��մ�&�M:@t��%Ns��%�$�b��:a�B[����pAh���J�֤��Cg�^9���Q���_ ���s�?% z�Nо�k��ts��^?䂃����-AJn�Ud����Gi��b}L�p{�rW�"r)���Q�&+g؝�7�T�� d\��$�L��>�C~[�8��!�����c�e�k����Q;��U���c�Y���q%���S���;���桪~(��3v����	I�J��%�z�X���6������ �$|V��#� \���ڌ�Ji�>DJ υ�4�ݚ�1��Hr.?s�}�M�)�UgLR�w,<=ݔ��������T��J��,���|a+�*�$���KL�d�P,�e#?e����6�$����{"�qUy�L;�/`�1�M�����QVϋ��}�� �'s����TRT��� r�+n����^���휼y����j����y�b�%��I�N�l��֣����$���'E��G���(]@h�)����L�1�Ha<>��+�-� 8'��K���J��)�f~�\fy�e%u }���$�>�Iܡ��(������sLأBc2����A���L��M�PI�����U��1��\[	�,��)ᤂ<����՗�/dEL�A�\��c.�\K��$P�.�����=9�7�X�4 �~}�e� �?�B6~@�7����'���*C%�&��2�jf��`C�Ӽ���0�����h��)���n��Wf�˵ꤥߨ�������ø(�ڦ���R��I.8N묃�y�EW�
��9H���[���S��Îus�S�/��������dz�#�������~��Ϊ�3W����	uמw ���X���"̡��+���0έBl���gh#���ח`c2p��r������7)�\i^G�0{ ��5�:�ErM�_����?2�6�n��7_������,���p�'����p��G�� �b@L��R+���������ϊ0�ՌH7F�̀�!�5��A�
���%�vo|��*KREC|d25�LR"Y���%|zo��{X�����a��[c�.#�X��g޸�����{�I�*��te0w����gH�J�91I�,��nQ5M2a�����h�0��\�b�Eڨ�^�n^�
#.a��uωQ���tԆl&m�?y��x�3)���]x�m�G2�H=aA�Vo�P|���� qm�h6�����	�x`k�~G�a�� #��3�M����Z��#�x��=9��`.U+M_�� җ���9�K���
�L��v��ᦎ�6��N�6��J;]�,_�A�٩7��J�A#���+M90Ɩ�)�$��~�H��i�[_rh�Ḋ �+?��7� ^�{�ޤ�\�|F�%1Ga�$�%т8��v�(���=g�>�O����D��>���?eF@��t��U@�(�Z�8�u���EW��y�Ҥ���5Z�����C��@Zm�Ҫ]��Л��IX(=j����h�O���P�zڃ)�#d|�ӆ��_� >R&��-�ܴ��Ϳ�'�xsps*�T��M�CoOQ �]1�O��Ie�Z*�>b�4���O
s��k�ՎqC0
|�CG�L%F�a�����p�$b9,x�c'�5��b�v�>ťH߳�|�zC�LEȦ�8Lf�W���ͧ�F�o�g�s��pX���m�@Lh7sVBZ�o��	WL��X�bB�S��_X�����o��	-7�PP}��To��[� |��C�/���݇��c��rZ���ᣟ�b�M�����1�Č0h[���nCQ��3� �Li_�l�ڏ����
��#�l&c�"��[�<	��h�+��4�TTP/6�1Ϻa��_mL�N��,np�"��_S0��I:��/�����p�%�42�������N�<�S�D�P���0�DEz�_Hb�o 8�ǰ�I̘���U�+�d���m�a���}��PMΈg�9>�s����dk��D=v�{�xJ���^%��S�;}5
r�j��6U�G=���c����5�/�R}������Yf�E+_ ��ĽU=��MJ��Y#����� [ɍ��S��$�?���^b6�s�E�*p�q���2ٚ���6���s�Ȑ�Z
ƽ��4���B:���%�؆�Q��G�K�<z����x%s����w5��դ��g(o7��e��� b)OB�8�X�5�WBl�PHA0�|�HR��\��7Y�dY.?ٌ6 ���;�(�q�A��}�Q�ʄ���'*~1r�X4�)�Ց��۵��=�ͽf���T ��2�L�:?��	����,6P� �p%�?�FOo�s�?��]�H n��a�у�%����ݺ�~�X��� ��K��J��-��d���K��$��RJ�`nXV����2�U�gA�F'OD<�����l�_�s}���-ߟ��O�!
&鯄�k����Rx�ڱ/Qp��q�ޮ2�G����{�r6���L+�C�|��יs��]�tz���T~vg|]m��=�� I�~�(�?s�q��W*t~��DJopD}��g��66n�nr�GcbM��2�>��n�?��Z��%|q��� GL]��Pv���SUH��ӓ�}`�֦p�PM^=�r���k����a�w�3Mس��+�XG��/�ҝN���v���窒�ʫ�Xc.�����!l��
S��{�!��(��S&�"tO-�o�?X�2�� ���wj쥀<�s�9�]){�E6�uQLq�*@+ �y��¼�P����MIJ�x�̆���v��C�~w�l�6�D�m��
���ۼ8)���C�8����<�{>��n�������|����(4_=�ʪ�~�'����S�y����9]���U�!:���ߵX�te�:]'�1P2��~���sԎ�)×a:-�<�HFک����h�^�>PX2���n�Ҏ�9�C�Q��r r�|�|�
P��q�w/���%�:jۄm�UƷ�1=Y�M��*��_Yw�߽�V	�C<�#ܣ�[r�%ێ�AI,=],81q:��v�2wUeſz����%�b�P(�o�]̍JX��/����F���h��S�|*�R�"�z�Ĝ���M�{\��x�'���؊Ϩ2��a�=Zlz�U�U�����eOE����1�t/V#]i��'H�fqYnh��?��@]L�*�Nht���&��Nwo~�{Fl�1�%��:58L}��3���
�p_%�v�r嬬�T�q��&+������;�W�����h���ɦ�C'J�l�F=
o!s>)���н��\����gM��� �-e��W��N�RAf�u�+�[��g�����6`��	���EbBV�D�V���!�DΊ�Ja�
�Ƈ�˾�Ϙ�֟y�� )o�1�^K��a�p�+��#�n�d����rw��foQ"�=�'�c�Q�Q�42��|"��п���Z".�VB>k�$��8�n�U�����Qh����e�J;�[��)Z�hD���naю46J�E�͂�r4����:��8V��d"F� S�����{	u�T����q;:����O��3�3�`qQ�D�x����c�%[��I�u����]���AU%��\�ZC*�x]�E�3< $����#�Q�U��H��~jњaDHɇ���QM�L�u��4s�y�?���u7��������;��/�v����Ӑ�S�
��M�<�\�t"���;���X6CN��vV�-E�<B��é��O�|1�Dݎ�r�i��É�4�c�޿�st˜2�lO���4DQEZj=����]�.�:����v�\������瓬q�A�M�6��4u��h>a.$d���Z��D#�U����79���au��%���tA�݊F!ʖ�f�k���~����z���+,>۬���Pѿe�.�QHEC���j�5|�}f�;s�1�H=!�~��N�`[o�э��:��q�p2.��qE�Rs�����
M�jp��Ӛ��J��Sr$���Pa��m�͸D���zN�h����LwL�KK�"\��[aV��:H�E�2��;��΅�0�Բ�Yc��n��U�3�g��ڤ�5,5���n�
�Q�{��~�e�U_�+�%�-��������NH1�W��~��^�<��:��v�^����d
��������.����W�����`_0��n���r$��g�ٮ]ys�KE��hJ��kn���=���r�D"�x����AY�t(o�77Hw����>BN���-�.Y��$|c�$�ht��Xtњ�=���q|�߲�?@U>��V�7�tP���+�x�gZ<�yK&��p�함N�⼇�A�0B]�
Sl�R(��;w����I����+�����8�,o�7�o1����#�n�V�b�!Gt�iJܣy9�㚫�;�-�5APq�j�6�I�z�4Y�:_��ǭ���k�����'O$�Ы��Ft��������!2����Nͫ��|q��i����	cc��o��Рp� ���P8�g��S�N�������gB��"q��<�i0�C]��j
(X_&��y̴���| �m��ފU���D��*�"�a��k��{�gf�����2TaX��]���S�Zr�P�y>{U��[����A� �-];?�m9�N� ���ަ;���P�L�0&%��ڊ0����IC	�v iF�)�=�����o��Gb����ؕ*Qg�|�9��-��_��DX%�:��x�<���o����w�l�5��0����h��|u�W��!zY�4[�^�~R8ٌL�C@no�#V�!^H�e�آsE�� �#�3f��p�����Y�I9?����&>+b��\�y�vl���_�3L��,�l�vt���0��z�c&E��g9H�T^40+�vrs���AG��&fp�1��]�sp�+���,C.���𚤯���?[J����si�_Пh�i��!1�ٳ��?I��:[
e9zi'�:q�����i�='E�%n  �t�Z����kp$&�3����h7���y�l�	�^m��'�b��+���]�L�!	�e��%v��ɤ���n��kt������_�s�J��0�ӌ*� ��bJ�fYØ�g�8��~�w&OJ�2ˍ��o�����
6]^��/A��!��n��YӤE���#��'�*g%?�̾���	��r;hd��/���� Ϊ�
��tkvW�P��GNSo 5�~�uQ����;t����-�'J�AOEhP��G�Ʒ ��`)�73�3��h�=�AJ�S���#(a��qQ`�X/��3%���{�.dM�6��<~�7Vw�����/p�Þ]ӣyp�>���������	�0]���h8�Ȋ�)R�8}�]�|;Ш��	.�@��Fz��L[���g@�7p��1� {�G���;��~�W�Oz�?0�(����I���h� sX_��"o����)a�~XOi�{�DN�h�[T�"�k�OP��y�H�/59������>C/&����p�D
oV���>��>���U�x�G���E��E�� �1�~7`w�I���NÀ��B[��֝R�$a�S�tV�!�{�[�%��[�6�*BG�ܾ���)��x��3B��Y�/M�/l�nC���U㊢�Zq�}ЕR�9��}w�<'6���v���~��4����)5+=�"��ڐ��x£��6�����\:�F����Q������ �%hc	y��Zs �+�_�!�3�v��Y|�j�3u���4�|��(��Wn�hW?Tg�w�f@ڸ�R\�34�:C�겿����srhA=�1x���UݫS��[��p�]`��v�M_(N��v`Q��>���,�+��f��|do�~n�BwE���.UJ��Â|Emz��	_e�=��> ��7Sx8z��4�w��L+��_���p��?��8X�d��W%;o�BZͪҟ;2(���$HN����_g�i���,�
�+�=β�5�kc�}����B۔�OM�u�����`VH}�k����;;.<��n�  �g��w8�<k��h�U�-��5t�-*K2䵪��%7Qa5���@��ZS�wC���e� � ��'T�(I��j��R�b:\,#
�0;�O���@�W�.1�.�)M�)����W�������G�Z�"�G�m;�k��(9÷��{�J��u4&�	hRk��.�B��8�on�(����)@m%HXh��^l��v�w�����9���UDϙ�W�������) ���5���'n�Y+���1uw1K�CU��b���hq���d�	��L�P6��^s}]�m�%���'#���~Q�#���T�e~��V��J=Ul|k�z��B��������@�<8^t0:��Yi��KU��7�&m����M�W��ts���!'W}��N�Y5hɕ�GЬy�ݵ���xN�������~%%��J`<(�=oFJ��8\UN��**�L��]̀TuJ�����	��?�x�p�<Ƭ��]�ңL����E�x�@�,�E��rF��]K?8\�p��j0��l��K�Z�l��P?�:pXq�v�7����Fi��8�E���q�c�"��q�3@ՓAԋ���O�*��8�"f	����R�\�.�ã��11������9$����9s��o��ߝ�Z��u;d��{5߇!�&)U�Yc9������U��ëG������Ρ
Na'B)���@\�����t�S~tM ��Z���Bl���l0D4�CL�u� �ًC�ayk挷HW�$�Cr�r�\��Zfgm�-�*��i1���X��������
ً��9����_dx5\n�w�䴦G���LR�9�O��Ѧ�`��ňf�������Y�EYډ�l�V�Y��ml5�=������`{S��9��æ�����@r���f>�����wQt]��ѩq��@�v�3l���H���d28\V��XrX:l��+ބ���/�HH�r>Ñ��n�2�/$�C��j*0*�Ә1ϟ�S���p8�'&���:�	z34=.�4�9b�->�!� {>N���w?�*R"��8�����@;���?:��ݧ@ 0��6���#t=b-���5�m/�&���@SfT����	����%^��}����8��YL�ld�W#�Ё-���A'yH�ʂ�vݑ���7xx?%���25u�*[?�>
sY�t��Z�������)ʩ�װ����p�!���ѷ����g�1�LW;꾔�uh���Z^�et�/�c��K��]��ð#\�����kڂ���j����X�s߯f�!
h���l���}�4z��h4�ǝ���S�z�ө�s�_ΪO�Kq�����i��F��֨��=�!�FkV��nx��*���*7r���lp�di"p!tw�]8��>BV�!:xg�6��z�q����Kj�(�����CH�:�~����?�|��c��`�(�Ø��l���!=����ۇ�	2�iD>�ֳ���í�.�R�[
��)a@ѭ���|�I�
G�%+���	��R�W��m�ztH_�Cz�bM����F{j%%č�N�e���(1!�%�5^��k<�F���׉���vI��O��k]��ԘZr-��`,�}��Y��3�x/`��&3�63��f�P�����xlY0�VbO�ɝ���UcP|�X��sU1�Zo�ϖB��H�ϒ=йUne��;)RI1���,?�����X'�Q-�KI��)O0^���4
���������]�P@�o��;0fy�5J.M���6�$`6��>����"ȥ���|�$�h�PM��9˃������E]�\��j�
qA t��Ͻ)�X6���,�Y��^�I���>��ZXdI�d�Qo	<�x�r/�*��د�П��_����1���>����z�u�kO4�jI=G8|K�Sc�7 P
]>���M�C@nZ�df=�H���d��7�7�c�L����/��'o� ���*`2�2c�q���.�^\�1���'�@��?��;��2�\9��ZE�+�$`�gơ:F�6�7[����WJ���q1R�\ɚ�>כ�1o�i�u|��%qS����9�8f=~��6��;J�d\;��ȟE��A/��Zh��hD1�S�p2F�~�T<�Դߥᚻ��T�Cќ�'�hTBt5h��V�?N__�^�1��'����jnց��3� [�?�8����C��͋6xڊ�H1�}����j?S�^U���N܉bM,.{&�{�!�ر��9�e0���%\�A["�l�����X�5�]F� yx5a���6R�
}�f}2��r@�t{��`֎��
�);������>������TcQ�]A�R�*�'7<*A��������|[��Jq�o�8�*�(WF6v�rr�>�Q0�i���O7��ζ�}�/0����)�m�k���L��\�1���w�Fr!7���ԃ
���,��F�0��.����[wɜ�S��%)>t�~E��J1u��n�d�TP��g�YSxD���8 ;,H��ĺ�sإ/�>�0u��I'�c����"<&��/�C9+Rm�y(K��u%�@� �4a�F2jf�h��Wr���Vȋ����j$�%y�ײ� iɝ���Ò5|0�TNn���m��'W
C�,�4���B�W8vV������}+�H�f��̓|�KKU�ej����G��r�o�4��64����#I���g\���z8ES��aX�.)� �1���CO4Z�Q��:��z*ͻ��RvF��^+=+�(���֗�@�����4f[��
K]D�F�<�nl u��_���t ����vd���[R��&��}��R	ݏ���a����R���}���bF���{�v)+�,W�d!��еt��#p=������@�5F�z���E�R�(? �k��0��`<�jJj��n0.��!�j����Rr���ӌ_��4e6��p&X�/s�q-��<cK���vE�����Ƌ�j  �ׯ[�!5>) =�>-L��(!��b�M��k�Lw���b���E�CO.RF�Ng������hQZ�zV7IȞ���q�;��v�
��*^=0�S���P�����;6-�S:i	�r�)��T�l2۸�Ld�w�8�g�!���dMLଭbb���QU���D[N9����>����ˇ$�*�-�3@Ǻ|C|
��|hY���K&q��>�i��;�4�G����x�gw[lwW�~�!,�<&��"��6��3nN��E��V�W�M��X��#"A�L3!d������"���I���f����!�����&w؃��X����5�qk���B��ڷi��l���.�ft:�U�q���EIecQ���4�8��>>�����9��[��xDu�A�a��*���e D��&	�@���|��qݟ8�ƝH��x��.i��a�f���K�eAN����]��L��=�W�O�σ���Κ���Ѻ��1O"�2�n�� ���X#�ٳ����ˑd��)�{:����,�d�t�ܿ�v�@��tM0b�!����.KT��=V� "�b'l�\�����wP7���fJ5+}W7�zX��,�/��~/��ߤr���>U�R\��y��_]��g�5��I�h:r ��P���؎����v���<:p��`i:zV�L:%'����2��J�6^�R��c#�=�	�`=p��ܘ�m���b"zY0ʃ� -j��J�F�.��H̚��������]��ޤ�N� ]<?y䃓^˗~LF�!j����{��$屩�K����(ȨO��}Z�;-IO�"i4�?4�^͂M�/�U`��7Y��Sn��C�bs�h[wS���?��y��45�x�1�B��w+e��Tz�rq�d����<�s�~J�xT�9Ń�"����M���KTɂd�g�/�g�h@o� ���֘��-n��
Tv����R��7��1]��~]��h��OB�y�d*�y��p7Ɗc���'�\e��q��bha��B�;K>'�rM�XS�4�)Y)V�ݯ\=+7�eV�	~��� ,E�j�A�5�7H_b~��n��<K%7ФZ�X��U2p��S9�@�]���B[�����2f���C�v b�i����c����,]W�a�:兿�³��̞�Ӥ.��c����/⼱��
W��
*�B�Ϋ;F-Ӈ�׍�����׷�{�s>S��ǃ���Y�|�MЅ��l+�-����LU�
��62���
�A��}f@���"@&O��w�A����|��?j�((�⫙喏g������l��k���)"o�	p����~]b�����8@��Z�1f���Ž��3U&��n{w�$�)q�z'�\$���uYH��;�����9�����Qn@P+j��v&Ӎn���*nbH��ɰ�j���
��m��VA$�h9k>}�[���>q`qu|�
����sy?� ��m[�PLRhD�٬c%�A�\e��Z6tz֛b%X��E�e��/�g�����6q΄�Y�mB˂��ʜ�I&QȦS��5W��o�5�4f��0�������1'h;ƎC|��N�D���`͆0�Y�e��|������7n� \�!!y�B���h���?J4,S�>+9�X�j� ��W�DַQ�\���������a�sJ̳��
��A0�ŝzZ�n�+��;r�at� ��x|��8�
��LZX0R$��spV8��KB��0�9t��`���@�M����s����z��v�y�h�.?�R�'9��˂`��_ӈD�����[z:o�m2�P�sJze�U�`�
���ǭ�ߙ��䚦$P�����AP�b���(��g"db�}���BT/���{sd�H����И89"G�y1@�#�,�����\��PL�=O$�ܯ|��ZDh�+40��NK_f��q�h�v�%"r3����(R�!JՂ2:	���b��yx��jՐ.��1���O��|D	M�],�*�\k�W����xr�RQ�S�e=�R����فHoAO}��vh���.Lͧ�:ҁ��<?��\�V�+����g_�E��a�W�i�6o���k��(�BK��6>���,��@��R�d6�B,����Q:A�zm���,��뺄�IoL��f���7�ޠ�{c���V'u΀|�kWR%kY��X�-��\�<	��ܵ�^����J�K��Ɲ E��w[}�Ϩ���(��)G ��dcKy��$t�d��}��G`a%n��I.=�
��u"��b�~�F�d�@�Ra�&k��<4�4�n��z@�/�j�U^xÒ��X�T��ly ���.v�$׽=�ӓ��T��(A��d��6+Mx7i;����Oк��u�֙��~p%XCM�Z�q���l�i�l������/���q4o�9�S_*&����O�����;�{a��.���Q�%_�n�5��E��H�P,^����l���t��LuBjHAD�6��ҳs{I���|�QC>�t�e/���ѱ������;�S�\�u�Ȯ��O�`@�we���G_��2z�\�54�`3J�a[����:���Bz��qRC��q�Qb���D�]v%QYdO�,���_�t�ְ{F,��KÃ��M��
/�1$�Fyh�L*�|�RZ�ܶ����Nu�L�,{��z�R����i���^��9i=8|���D.�B�4��T�N��!\���ۚ�/�d��blϷl�pl\&�%O�1%�V����P��t<9t�阛�yz[��SmP�"'2��^S�FB�J�]����7ږ�&�vF&�� ��!вː돩Ɩ�4�L��Vq���������m(�բyR�N����8��g��m��Н��V�b��" �����2o�!�iE�ݥe��I�e�K�����ӽ��zھ�à�+s#	[��IƔ��魖H,��3�g��?'�!�KM�a|ɉ��~�#J��G��ӣ�[��p+)1�c=�3	�������L���;����<��)#q��F�����гk�W�¢�p·k�N���/'�g�"�Zt�nGYLl$��Cܧ�<#�rv� �LS`�Xh�+;�7-��B�b�+-�yX�\e��0?G��K'�������"ǖv�%�ЋGp>��Nv�3�G^�K�P�ţx���H�?�֢�?�ٰ\�E?�ِ1@���K�%�"pgf��q)���%�^��@T���a�i�iyN�[�vʋک8TP��فY8P��̥�|P躈�m�Qx%8��s����͝��,��ǳv��0�;�B6��H���P-�Q�:� p�t=�<tEU�������f�+FG�j�B���哙�7wlϝ��(}�H��2�	�U �æ� ���7/�%͸����6�Z��A��)��چ]w���׷�'�&@�%��V�uI��^�,��Oo!W!'&�\��w����Z�O��!����_PI&R�~+�EY�։�9Nłý�'�v�i��]�v�>qvY��|TY�c�iS���������� mOR]�Φ�B)�7�h���;!�[�w���8a��YCy)���{���h��H=/ �|��x�Hs��>kE�*��8=6G�5���+�Fcz�w�^����Q"�\ĸ�Y�Cu(�I�����U�4x\����bB��9"�Ԃ��	1������Xo�PF�-�T5nf�{�@����������ܼ���O�\�odF�� _i���|` K� 5qË�ר`���H0�_�����j��c�0�k~��(S�}�10J����y0�z%0�L8�8b��?5�ѣ���[��ds�H*7�z��N�^��J=�d�9A�sv�J�y!L�]��l�{p��%�I}�	�~�J���*��R����/kR�F��&�Ƃ�Lܞ�$��G�C�+8k�iUi�R�c$6I��0�t%� ���ڗ~��?�z7Fk���Y��$�Q�L��9i�YkT����0��ךSuB�M!a���F|�K���#u��4F�(I���1c�C��'71ͳ�*�w�$�!Q�8���B�"�Ӆ��EddR�gE��.�S�(q����:.W�D�鞃���T`�>��8�u`%.v���Bq�TR�R��T0�\� ��ݼ+�I�nv'��FW���j�}.{���'����M�vLJ��[_�v�����1�:6O�z�3q����	��pg�����TO�K��7�(F�UϮ-I��\L�ɲ,�P2��?�NG��DI��)�v8���V.��v�ת�����^e���cӍ�[
�P�.ׯ����cQ;<�< zw�rJϽ1YX�vg�<F]Y,�o�}�j!�{S�B�#V�f2�,EocpTڕ��Ys�n}��D���+�kJ]D��/�:o�&��U���/2<��91��Ӕd�������X ��(�QJ{�f_��z�9�I��	���ټ�^�c�	l���'nn�/���A�d�ն�$�R��sT�1	I�~�b�"��&ۣ��,C���	l̥�y�j��W�{��j�'r�{A�s��u��NG��
qh���]��7�S�\��>���B�+��Čֹ9%;�Qh6p�^��e�d��0Uq�iV�c�^�� ��-�-1�&��\*cg��^<J[n������F(8�UN�hd�+�(»՟Y`��>/�)��d���,��b�t���#��� �5�'��8y���d4��j^�Ar�y��\خ(�S5)�V*469z��2��%���}��`t�h�%'p.^vS8��e��a�Tϛk���u�}�ׂ�p���ca��}�
�)�Gp�����h`�8l�ƙ{����m`F_��x�>�"M��4��s��� ������o�n��[J�ǹ��F��c>��M�� L 9n����@�V���J�~�=W�RcRu:�����'��U*��Qh��}e
N���c���ɰ7,0�(�o'(�b�h	C������h�m"t��,�L�MK�q/�D{l�Y᪄�h�Hzmi����<n��g��
����L�4|qb�`C�{�-�(b�K|�P+�p�n�94�ع��	�m��L2��QP����t�XdQu�`�B2��r�?L���c�U��-���^P
G���.Ni9<_��w���L�̃ԭ����2�����w�K� ު��I�=!y�^F\����WÞ5�9Qq�:��[]k���#9<���(�{�B7�����k��jQ��bH�+u��x�^}gaK�?ح826R�{�^��y6�\$_�"�.���X��E�Lf�L:p� ���g�
�5XI9
pS����d�ގ�ςP��c#�k :�H�#y��4�s��^�+��T�g�t2�Ŏx��g6\��F�[��5��
['q,�f�V@	��l��f|����x���P��{�ʴ�mb<!69��xnG/$5�`Z~+y�5yAG����o�.{��������:뉒�h�.��U���;�ʬ�"8;[�^$�^��U���.�a
5k�C��KH��wI�7�׮�ζ�ez��dh�+���6��%��8Q��",��v|��c�.`���[k���X�J����Kf/��/8��!$��;���5���*}
�4Q��8�����G��� ���!���r
yC)"H�� -��[��:꧘B�6��R�����T�Q��c+44��ą�G$�;Y�k�N�x���X2!��2�	��H����C(=�Ҿ����`m�.T.��\ݭF��Ag�H�	6 �6�(���K��F�Ȋ�ZV�C/�XQW�t�Ӹ���+�g���b�DP�g[g�!� F#��;_�Rb�}ծ�l��'��Fm�5�����j_hZ.Da�׊R�y���νH��3�xJ@�8��liDLo���K��R��\>*�Y�!jnȥU���[.oRH�0��d�z.V��=�X�ݼ|V�=��%��x�Dv��j�C�����f�g�����%�L$�}ARwH���P�v�n��~\�E$��8Kg1/�{��	g��������t�N���K��e�F��
e�����A� F+T���A��O�d6��fDv��x�p��*�����r��{
�]�v�{�3��=Y�;�����(�πSF�
�f..��h��д�J�m7|�rG��-×'�:��_��NB�W}��`��2��.�F�>X���"��lEOo-����wƠ!�aN��M�SN�K��'�˃���"o�z��>�t�d��0�T8�s��������}o }Lֈ)���1p�z*-6ݭ*J���E_=�td�u�\�?�Q���U�U{3�`h6�����&�B#?
 =�;����n
�����,�6��������T�r�b�
N�ۅ�;5�c��oiӋ�3���n�
/�dŋ�ĀdxN��D�L�6J,�����B��pl���bb��қܲ�L��'#B�b&�&�~t	e^��8bd�e��<tVMr�z{ˊ� G��#Ƈo��]��W3+�D���YΚ�\Y�@��LxL�_���P}E�2{�Raˈ���MzC��?�߱�o������U�+T<�Ǜ��ە��C�Y+��A� x˸/��w"����fM������l8M��b�Sd�2��01~�aP�@Q��UR�ABëMX�~����6� ��)�uUD��w#��~�mA/�r�xō���ڐ�oDz��j�B����X��(��v��o�1�/"�C�l.1~it��������Ӓ�����-��Eq[�N�q�U�
��u�V�H�c�����u��`�+��G�H�$.2H�M͂[�f�~�V;c֪��/IC���u�L�F����4�I��B�34�E/� ���p_=�� ��
�����^�:�W�V��۶b��]xJ�#}g���Ze��|�����%��ܸ�?��h��y��SW7�����#�E�j�T�9��#C-�k����9e/�_R[<�i=���V�#�0*��7�G�m4f�M�k�-���[�RԀJoC����p��̮Ga������gY�B{�=��赾�U�_8�ԉ�ɛ��z|	R��u�`���^AM��u�D�/����h����@���R�a3�I�V�ѭ�c����wN���U�,�Y��!�NdvJ8���}/�U�N� H��7X�t�l֡E�8\�i�S�}��w=7��F|w�e�S"V�##�N�����cH�S(I�#^�[�]��V@#�w��
�6W��z�P<�z���?Zm�
�+�,T_=�a�dܿ�|��v����ך��H,�s�O��cg̩EN�P`#�OD�H^q"+�eO�������5�<B���X��D-(�������~S�]WBY�ó&5��aߩ�<=o��<rz����-�����{����`'P��V"K������
�AA�Y�Zx׉d��*�����J�8�5����F��Z���W��"��Cn��Gz�Y��|7�����к	"xi����Af�@�<���Q����y�i��}?g��c��$�K[�E~2�hr鑡{����Ig�~ЏVG���rǞ�O��;�Fj�-xe��ϟ[�Ȱ&�*C��Ļ�]3�B��5���kw�0�e�b���|�����{���u�A�V8���uqǍ ���~7䩖���bH��/�Ė3��2�`��yf4E��w��j�}1��c�&E���X��!��c"�6
v��="em釤�r���%�H`�Ⱦ-bq^����T��:y�E�>���j\�Nrc �T����3�M@Ҝ�4s��B���/��<&�a����U�D%A��F^o�/���(I�=��K��n�IMJ��T8�`o�ĉ:��՘��N�&ӮB|܂�'�B%�[n�z��x`��gOn�
;:s��a�6:nx=��8�֨6���$��}j.�����h�3��&k䱫�ZS��IР#�P[��[�b`~��N����@Su��[�����-�#�$�C�� ��w���Ƀi�϶�B�)=��+����E���k��㠚H��nK=��8m2�@���coȯ�u����T��$O k�I0t���]���|�=������������~�;���(?7�?�guJ���2j���-.'�Ԉ��en�1wz��
����hG��?R\�)VN g�H��J� &�����S�����t��O
���ʘ�ч�P.�j���=���OE�ӬP飝G)띻%E_�(h	�侇�4��y��.o�.u�H@��$�k܍�\��E����Ot =4x2��%s��������2��n=�4o����A�eј}����sT9v�`#_��ȭr����:\�ͱ]��<��6�xv�a��́��2�:����K��c��b�<�B��e�k�أ3�@������d����(�n��T���	�=���b�"�p���˅�����MCA�����d��l�?x�ה�rr7�P:f��̏_��4�}���V�����5lUX
�􎲦���i��S�^�@�h�m�X�y8��fS,��f���<N�ڙ��j5C�	�9_��|�x�@R(�
4'��r��U��kͥ�liYբb�i�.��4B�}`���3�8ŗ�W��w��p����"��	�4R#BI������bC�e����,�ɍH���I}W�����B��(�5<&�> ��n�ͣ�g�BJ�ei��q���y��߲����0>"�B�%���T��&{C�ر�.X0�c���s5߹�U1x�W�'�˄̉����u�b��9(��2�I��U;N��<�R�b���H����vڛ�py�C�?Ie̓��U�ny��;�S���6�9�VT�hjYS�}�PJ2������4��͟bywH�V�泣��+S8�b��@�f"�[TT@��\F)�=���xS���� 6�ʺ���K���eߨ0����e�A�H��k1#�	�n�bT��n~��<S����wrJ��pUW,�ݨȲh��fd�$Nbn�����?C"��|�k�<��ɲZ���9~:����3�w��V6��-c�Y�O�:s =�Qn�5��������w��Ҡ;kHrR>����X�r<E����d�tx�\!��0F,������N�#c���(=���31h���]�\�eY�t/��(�jz`�>�u��U�L���-�OL��{hj�"9'�4\�rR�5���Lݨ��9=v9��v|��3_��0�`4�I�O׮�gk��L-��[��x?b�h�U
9mI���4ks_%d�r��s?��mp�y�	B��r����v,��׼1�������(�?���NѤ6�X��m��Uq���8Ѐ3��PO:�S;.k"	S�[~�������1�I0�7��P%��l��kd
���&@����l�B{��q�cV�J�lC{G��+�:?h���G>H�!l�%�I`�E�T_��ۏ�K,IT���8��?j�LTM��Zo��F:%9�>m�7�֬���� �`S���j�3B!"(�Ͻm^��
�x=�sn������|���S��q���Ά�-4�����'�ݴ�^==Q�Q�e�m���t#҂i6��W�������%�� ��*DN7�AT~b|W}�{��R�	e*�9F7^f�Kcw�m��t�?ſ��_}`Qa |����:#�N�c�Z�dIn�FрC��Uz��� lQ+\f2s��Sr78t�$YYu�FF��-' ��W��W%�n�6�W�6q��K."����QTt�#����<,�J��>1TG_����ș��wۋ�o��V<:!�Q۟�t3�?4�?:�j�8����(��]pZ u�6���&�e�S(r5�pN� ��A���RT�;� �;��A�Q�L����˵eW����a��.�s	��/J����*�XoS��O¤��E��g��N���ϔ��3�3��<�KTP�������	h�wS#�x4c��Ԓ�OA�T�X�=c�jC2��-�/��坾i�қmM�B�0�"O�,N�����j��|� �̦jJ�#�
�R��T�:�ˀѫ��V����6P���ទ��_��{:D�PҤ�o�߀� ���� |�?��z`{�ҏ�{�w!�ot!	���)��-�"���|M��Ԯ��F���)cN��~]��"�	7��Y�Jv�j܏��3�Hp�����b��E�X�%�{��1��
���,�V��_69��>�m:���I���n��Afϖa�9�ﳐ�|E��V]{�3l�*Nί��C�4����uFi�KH,'ae%wT:�(d|��*G{����o�h�x���kp�`�i.i� �����}��*���øz�h�%�J��/��S9"�[W"��/��@�f���x8��w�P��������dS��WM$5��'dխ!kۂDbR�y��o0��sa6�d��M�r�r�h��i�ܸHSݡ8Z|a�T�X�}d|ݚ~_F��ps�zp����0>Ll���\�!L�� �l�����|��ҍ�b��{��,�M�=�y��J$��O܅�J���M��{�\m(뜈���(Ow�~v�`,�Pݓ�������S
+?T���Hcm��I�>0�O�Uu�����nѭ����clx��:�I(F]Sg]uWc�d;��<H���7���m��#�[`���&��:@	 ;P�����l_���0۰>ԓH3�]٢��V�d�:���Ϭ,󽎟�DR�K��C�pdb��X~)%9���H���R��E!ц���ܕm����Y����4��42�pA_�C׸7K0�Xs�M\AK�g�h�Ƌ��¡����p�Iy�#��?�
_�6��
($�p��j%3x]s�O2���9�ŀR=x�n��~�.}�q�J?��ٖ��4���b�+�w�_~�y������m��`.{V���"'�F���V�E9�f/�T&��X���˱�E��^Pzܬ���?���e��s��B�Y��
�r 4;E��	�tt��^+��e�θ��J��cP����-d{�('}k-����YqTH,Zs�2�0A�R֧>u�l�4xVm/�gQ����s݈�Z��Z]�P�'�_��UF��ď:�	����J�5jS��׫���u9l�F��N�U	��2����5���PQ��1��|=^�!i�l���nV)���}M��dH��:��u�V��I�'�O��g���7H,+�E��|u�m��t	��3�,��S���C]wM���G����4��떥lxLTG��/'�5lfH|Hp�OqK��BwGQ��;Aa�A���x@W8*W*�knsI�����z�x�4�ڡ�VMd�c��_�+Y����Ikdg���T�s�!�T���g�EA��Q#|�cY���IhUJ2�n�C��%�<�\yh"�W|�N��!r3�\������9�
#C�R?�X�]]O3b����C�a/V0i��~��c7���ϼFݝ6�e��m���E>yG2Rc���X0��k��>_5Ԉ���Qn4pwLm��=}B�/q���:|^y�O� ��7Cح��р3�[�)�И���=�^P��?�.<G�(rlc��9�E�?[�e��w��~�g�^+G����z���p�,J�r5�k��Tb<_�Tf�v����P��l��EB���[�j����]����}ʻ���V�A�h}�q�����Q���q�_Cny���^�����x��|�,��˯�h5�1��R�I�M��-��dO�����);��4�^&�B`)
���P�(3��\!.�:�:>�0�h�00����m�h۾>���.|/re���M���{+����qOs���10��)��?SPs:��.&]�
���`<Yʆ��O�q�_�C���9�LƜB>�z�b��f��@�"�V/��A��~6��(>����x϶��U2��M�w�F�?nvZWjs��!+�i�QáN�KƲhq�>��7�,trqO��un׫g����m��9��X6��A՝�<�$M2�%7-^@��f�VM=$#��0aP��.���6��qg�u�Cb�l���a���b�ٍ] �b.�	�sn�R��~��	�RhC�<B�����e�����z����q���*>R���#E��5����n���{���Z�c�r��=�غ���Fe>�M[�@���k��K]�Y�N$V�8kvF��R
����2� ?˥B��'8���D��)��d�#�����.��j������|]�D�i�'���z��w������К��iB��6��Hr���L��/����VeQ��`�j��N@},k)������_��Q�,1�4ߔ"5���̧�K-�|����ȵ�Ms��aÙ�p��So�b�}�C��T�iͷ��X4���o�¬*�ΛKs���:���B;b+VH&�4�bvZ���)5��?7��:P���Rn�J�h��lƹ�g��v����H6���,v�ݘ�d�V�`�Śg5,#�ۃ��?2��
�|t���	L��OP�v�&�ߴkQ|��*��c��g;���e�=][�c94?����F
���r��ڷeA��?�4�+ث�@tH%rwb�:(b&�}f%v��K�*tBɪ�����׬T�ˮ%C�҉�b�Y8���:��W�
��ZL�"e\</f��m�3�D�-I���Xt)��1��� +Ϟ�LU��́���=4g��4m�u�f,'Zҩ'�����8�r��$唳��~"��E�yl��	�˩��1|6�t�����ɜA�2��
�}pWhf�,�>�MJfnL"�pI�d�9"?5��)~(M]���O�+Kҹ��J+P�k�\\���z\�h�ES�!�Gw����K�+��]�i��NOxb>�)�l�I3\͵���A�B<#�P쯛�J��y��M) �-͇��3wQQ՜�G�s�V��6Kԇ��Fݰoy�Z{S��7�Q�d3/x���$#x;H�s7�L5(�ۊi��ͳ�3�K$��p?�Wj��n�`4cE+�egxI9@{#J��m>��v  ���ǜP�g��	����	�=C$��$Ofe��=�)N+���!��d���z�a��J�L��]�"���C�/m�'�`8�oW�ǡ�yT����/�a#����d��H�jYG[;����o�{����xxh4� �{���+�~h4�f'�A���x�*��rX��6j�������@�f�5�P����3� �:�L%.(��2=�U�N@U%��Y����zaX�6�lBd:���j�R�U�a@A5�5�zY�&��lI���k���/�켎Kq�.�6��1�U����߷��U*�+ۼ/z�K�2��q^�2�{�� �3�{��v��w�R�L���qB,���E �o��|���}�"*��n���N��p*�.2E����|�6dT'5^���b�Z��1h`��������ȿ9�}\�L���8�R�\���K�����q"T�j\�њl��h/zeڂEO����ore`�Х<���Vh-'۠���۠�ֈ��o[ů.aN޴�B7����a�]r�qN���Dc�Td��"h�^tx8�ɩ�=�gj��~����kA�fO��݃��A{���ԥ@��q���Ҿ��c6�\Q��R f�H�l�@N�E	 �����w���i\����F�晇;6��c��n�`�y����#}>̥-�W>�ih�9�J� psV�n��	ͻ{6ָ�|�;B��,��P]��r��r��%9�̋�~� �i�A餗��}iKFZ����o�l`G�����!h�w�!��MZ���`���d ��[N���s�̷_� ������~c��=��=c����|����j#��Wq2:>_M�9���I�2���S��1MoV��+�M��]}q�� zYR��v�v�����>�U2�Zf�Cb�']���">�\�5a�#�2$n}Դ���wD��9c��`:���%{U���H�U��	 $���t)Y�q��0t��IXŋ��"&f+������%[���GA���a���x�
���h�'W�7V���s��{?��R&AA1�c05��=9�S6��qE�V������4z�h��U:$ޱ�sF��:�f�f��Ĭ��zSpS��~o�<h`Q�!��"���ۃ� Q�D�@�`0[��h�(P4'/9mZ|#u�0��!��xDVT3�X����,�^��{�B���?��5��R\#�[T4d;��&2a�q�?4��T�U���!��:���0;�2%.�h�j�}ȱpOYn�#��ۭڍ3�<b
�SY��*���3v�V��țnK�0k9��ž� �9S\�3��N��"�|�˪9bʍq{ �X�1x0�hp�B�q��P��n��j��0�n���ɧ,�1Ab�z�RcX񲇑�(6�Pq[l�[��/�����=�
�)	��Ʒi?����Ԁ&P�P�[֜Ivw��i\�xr!�8j'8�����|w.�t�6A��ͱ?Nj�[�:C���"���|�t��ˡ�}�q�A��|�*���W�[J�]*Yb���"�z�R'�+��P1��>����{�����-#�CK���ZW�.�U�W�������-�WTn�$B��|��Z����6ɺ���g��?+'ΰ���w��/n������ں'��V>z�@�.$�\ ���L�Q|��'Lڨ�>#ތ=��������8i핢�ǜ��xO���k)_���R�F����*4p��Ix�[l"������l���}�v��_�5c���"QS��M�>�'k�Ӫ���Ea����u&/�t�Ute���{o�;�E4�C^wC��hJ�;�r�<~ ����N����~(�q�g���n��S�F���Dz�h<��P��"�P�Z�oO����w:�@��F��j��a�+��������[��y}�1{����]Le���&�P���f���;��ņ�����kM jU����T��չ���n�j�VE�|R*wtz��er��<L���7߶��_V��Vff<��;6�Ѿ�uP}��i�h��X�2��V�b���/	��Y����;�/:�GU��B-��/_�C&��S_�DJ���$@�=���8\*�����P�T@�����A��>O�p���17ʀm��Ϣ��Դ��d���a�y���ΈW;<�e�L��@]����_P��E6V��27�f/���k���w�u��8f@w4e����8�e=����������V.� uN�X$��s�O���h�� �e����2�%(�:3D-R	�iX=`�O�fqG&���E 9���܂�dU������k4Rvқ��	ܦ?�OQ[$��dIes���'�³{	�0���!��Or����^�kTg�ɀdܐ<�oq	�_�F̓U+�~�&�e�0f`�`M~W',�"!GYuLi��
£W<��`���v�1Fux׊�¦	�@���[�=�^k�w����H�:��K��I��W�V�J�����w/��p�e$#YL$�z
�q�l.(�/�ȵ�R����x��R���(�o�i3Rm�ģ�`e��(d;=@' �����`����F�^RI�)�#$̝�|[N=!��6�4�ȏ�PO��df�Ι�>��7��ۧ��>= \5]c���ƫAy�*����|�����O���ut����H��8==���c`��t��)O���A�Ϟ C�|eǃ�"���o��du'��zw��0�~mt!�37�/��=��<������v&�X�>�^	�\���Ȓ�l0���K��ù���ﭙ
��y:~&���ӟ��a��=d��-�I��,y���`n�zR��~m:m"-P��JpE���٘3��l������Q��MV��R+�.���+�ZT�L����HC��n+d2�����N,�ߟ4T=�}���
�1�n 
�E�n��r�ȿ���S8�(�х`�,G䟈^K=�KX��dP�|b�2F�OEX�=$���Eu`�]�:ּ��);��;�,�}�Щ"��Ex��(߀�Y�����A�u�P�TjN����,�2�ů��o���2m���d�j�0C
�?����>�ҙ�sY��5&��X\�rˉٟ���j�M�[�� �M���3���%U�:�Bu�=���-)��}�r�ޜJo����`�o�Q��ٝ����4���ip/>;��0���h8��c��J Po�\2f�o7X:^��xc`�H��x>��ܙ*&
�EV�e%q��hc��<9���9!7��rN�@��3F�4Ǌ��:����u-U�����{`Q�k-:������%��ڵV4�B�L�`]����B�N~>0E�e���G.�2����%	{d����9��	��3f�� ���Tnħ���~��Mf���B���ʏ�-�l@)�丈4Q�:�R��ЕI�]8��M
�b�X�|�z
�Rm�M�`!+C����s�I�J�(����1�8���V�:`�b�����mr�M�=��gu�Z��,��p���y����k��m�����Y�ȩv�R|Β�юEc�W�Ό��"������	�R2a|��4D��-����M��_��
_a�����򥜪�����6��ӛ��c��l<v�
�D�QdMS޾���̸*
��1J���F�E�=�2�<ɞ��w��k{��=~�8`ݸ�@:�7Ymi�i�Bj�E�D��,.����i��5kH��=�~h_�=����B��A��T�M~8 �@�Th�kp��0\��g���	��`�aֆ����%x�5���T���g�q��~kiX��_}(�̛��h$��Ql�^jC��I�h踏a� � �X�չ�byQ�j h�Xt!��*���KE�|�8;?��!D��v�?�^r)�=�F�ܙ^�u�S6���.L���<���V����-�#ߖ����(���|?�|�#R\BOӦ�F��e�l�C���K��q�G�3MM7�QJ�O�/8�??T�i�6&9*i��{	���Z�֚�[_���1�)�vٴ����w�<q)8���l�� #m�\F177�Z�|�2y^�̧��$�&Q�a�h��67eu��d�0�2�Dyp�Kd�0��� �ס��[
�3�3R w���H�+nqj�E]Ē3TI�J�'/o�o� �b�$6���dv�h��wXy���R�tV�/�.��ms���Г�n^���}�Dee�r�m��_�A�I�k����᪪y�E��D�$�������8�k4�r���_:[Ll��˂e��2�1rH�/l���>(�|W�Ӆ���H�:�R��>-�#6�{�a��X��@���ʻ}]�\�v&:j�O������J�'1��w�ɹ���As�^���n$.�Ѣ�g���@�<�_�=ֈ�1;��V�o��i���෈�y��Ʌ�4��[6"-�E��z>�Y[5	`������6�,�Dp���_k�j��ȕ��8����j�VH�g��\j�L���o�������y�y�Ԃ;ؠ�*j�۰�D�=�p��Z���ȑF9OP:��v&9�����Ʈ�Qa�gp$�7����z��vD! ���Z�"�'�����6X�^Ѵ� ��?�qa��k�|�{��z�gh�o�÷�|!3�)���FN���i"�5�j @��Mh��*�8(�s��ֻy6�i�2��uU�����G��rY�J�M�cnғ�8m�"D�TR�m's�����v[�����m�o�XFȣ�nFO������s��ĥh��nO����Š%�����N������W���U7�1⺀Q���.M�wx�����|w�1�X�6���/Z�7TL���$�!�{�C̨I�T�3]�v�h�놙b�|�x�wU�%����&�T��@?}��7^J�M������X*�W��^ �cB��C'6�[�%�-���bz�z��`yc&R��ρ��-�Ƹi2j����ԽS�O�O�s��`6rM?�5g���Z�W[���*>���T�
��I�"h7��U�X0���aM	JXС�ƽQ� ��k�~��Rf ��
$�L�Cϯ+,�k�a�Q��<����[����M��\w��|m��'4�@�9Ed�K�$ŞR[��Bp���Ȏ;���S¬�r�wA�����0a3����z�ě�؞mi��P4��� �<@��_�)f��Al��$+Y��F�ͭ{;
z�'��tq�Q� VF���5jA�k�����;ҏ�����~�El����G���Dʃs�[��~:nW���{���W"\��7 ��і4Wa-X�Y�9L�rN�k��F�t���ix� n�<p���0�c��	,!UۥONK�3֏:�P@mԇ;(ao�)3W�A�%0-��>(�m�	>zD�7B�
�- R����c��p�2�*�vЫ��#�H���$#sl�-f��}�����n�%6���O�N2��3d��n�[�V9�7�s�W�����&[���̟q�a�pS<��c�����^2់R�{��&?�=	����֨z�m�l1l����+�Oi�N�㐛rB�\K5J���r~�Q1h~b��"�c������cԬj���$f"�z�H��~A���MX^9�_�U3u�n�U[E����mL�$w�NP fHq"J�F�x^{A~�n�W�3�����Du����D#Ñ��jnO�Y�J��+� ��&��UI��i.񢏝�=3��"��{,D,�6<�H|�T��� �;[����|�����0�%U�RR=�@�K���jջ-��&(5�B�;��/K�M!W��;����X��XyN���Q1�|�ܖ��lcE[�M�El��F�gs�/5������T��bJq�h�R�;��Q�T�l@���b���q��K'��=�Q��3w�,����u�@��h���b�4\!WP��AB�=��)��+�-����aܒ�mUU����֞D�ǝupC%��<V�V������0���*Mև�x��:2��n^��n9G�����)ޒp�ZW�N2�V	���R;�I2�i�Bw�2�)T쓦��|����=�Uo@�p�dU�嶾T��%A��78�K)���dх�.9&���|����z���-�сx�jޑ����}�i��
v4�詬V�x�%�:ڢ����^�vB��4�3�z�\ٽ�ɢL>�k�������Y�h�}kMSd��/��wX��w�U�r����s��o�A�Py6� =uFY�3�,�Q�.�O�#�:�ꐃ]��ן@��zI�@Q�oߖ�rB�6���5���J�BJI_W-[��m
0)�|!5����;�s�Y�(�%�$�Ă�v���R�r-Y��p'��W�y�y�L`��`�����-�����5g�Il��ȑ �����`X�Um_ԉ������
G:�x$��B���͓!2R�5���Up��E�O;�x"Hl�tc�1��(k��l6p���&	BQ�O�47�����q����j���w�8��R���7�K���ɍ�|&s����!������=��=�I�w�����;~����Wn���l�?{���%|0���;߹���"ۊ�Z�Ɂ?�b����
3�̄�>a�����%�rC�����X�2��fu�3����|�me��sZ�_��R�}�&
����Ҧ���y�׹�8�������x 1;U�P_��<�*(�˭����}I��6���{N�[9Wxx��.�|��=lE���X��b��0�ܞ������˃)���;�!A��j��wDT��q�Ǧ������>�s
�� 	�p�NrG�_ l��餷��7M�.�wt��cRmPV�����ށ2~���@��Z��G�^FOBGT�ϣ�y>ߞq�vqrAV�<�\�f�$k�(�E�M� J�W�J�5`L��Q%'��s!w�mQ!��G�|��ba�$=F]�&R�h��Q���mHP٥��U~�؎M�'n�f@����Ky�p:�<Ʊ;A���c&�t�V��T#RŔ�?�W
�Ko6�����/e#J-��4h�pwk܋�K�X�6�3���(KWC��_E�"���"~0J���@�4�]���I;���×.�a�#>�!,u�G���.��@���i;�u�w��
��{��(��f��Q��iN��a��<�I;��e�iy�c�����BT�"z��xs�@�[5�ݚ�Z�e|L�3��I<j�a�	�_�$H���f,<5r!%�U�H��%	I����]����	1���[0���I턡Z2�`��ʉ���}��!�� D �6}8I����g1�ps8�M���BS4�iH+������nl�������,c�:a�*ձ�쀊=�%hqA�l��/���1��.\m�&:z��������X�����i��Q�Ӝa�.��3,��c���g+����џ�5�o���ȋ֨+�g�fm�;d4Nn4B1�7{�#"[kK�O�{��u.����
QY�}$	���}�e�IN�u�}�9��F�]����h_�p>�]E��*��r�W��G���J�^�B��� x�8kZ�d��?�"I��, G�	v�v�j囍R�1pM@��6�(�`�ݨv0
?ۜ\��=�y��>��Q��R8��0<2�@P\{���!�l�f���٭����I̩=�!N�M�w:>w���7�\���L�h�u��\$��y���cJ�X3�E�6a���6�|7����y��P߳!ެV�6͠˧��.2F)+9.�5@B���?'S�G�e��LY�(o��XA�S2��	���bp��k��:&g����l�t�'�֐�@��#���--G���V<w��d��@D�����2���?�u��A�"Z1���8E� �,ޞ���Q�Z��8��G[ȭ�����3�w�I���7l���X��l�mX��\�Q�rN�+VZ�Z�R^������/�#�x���	"���3�P��&�6��=�9�C���E�%4	J|nD��ϸWrn�E�/���}����7���B�Xj�"�¥�.��4�
|]���0
k�:���ażZ��[���д	x��*`�z��u��KޖN18��&Î)�iq E߆m���\W3��U����L�6�� 8 l��=L@�K���<��Gd0�Ad��p�^d'@������U�K���Mr�X �c(��H���u>�Cc7�o�S���Ŋ&ܛ�M�)�ˎ���d�`�H��� �ǈE^︠$��W��� ������w�>^C�{��=W�F����c ��_F-�F���M�ue�0(�o8��\���G�&�Ze����创Wʂ���G�r�j�%�����Y�6��h�a�$���C��4Fg���uN���؞N5�n�--+����A(��<�>$�%�q"6�K���;R�~��QZ��SNi��|��9x�/�F��P@��y],T��M��=���y\1��U� ;��+�ad�r���S��r��R��J�R�I��8��ەV�E^�
���{I���c�j��¼�`��S��eEg�1|�P�u�,���/Ps�k�M@��5B#v���i�^��]�<}U�vB���C3��������+J@Gg�>�I�a��f=�1��5tO�-L��t��)T�Bc?{ʸj<�+g)���W}�If _��X�q,��_d���e~�n�� ų�>��V��+�hG�H;U���E�]�`���4�?|�ry$V&�L�b
6�����'J�K1i{��`��$]��7�S��W!ss+�<\n����M�SqT�YOO|�#̗�z;N�@���Ufc4�Ⱥ����_�⢅�(LE�m��RU�/xpZϺ�{ -6j�j$"Q�:W�6���O4���S�P���K�$�/]��1�!c�G�y�)��Zj`��҇���
�z��H�Ș�Xm{Ow];_��5-�~G&�����2Z^�*�J���񟪰�����!
�QȆ�,����G+Ǒ��̧��!A� �w6�a��V��7�+{>����a
m����jB�ɸr��v�6w��6T�i�Dhc.�7��l�1�<D�}0�ZI.�uo� Ŝi�w͏��pI奰B��&�6�r�W�2'J�GS��o!��d�џ��r�����I��ptJ�:���Y��P�P�(w�8Ò�C�)�S_�e4B���~3�
H9�.βe��6`��U&���r�w."���9���<k�(7�E>qA��49q���j����Q���H6�2�r1�p�G5���ǔi���ԁv��i��@g�M�ym<��@����mR��Q0�[�BV���%�:���	��$}1,��v 	[A-HQ�v�q��vVL�j������J�J�]����*C�I��X*����ڛI�c��Ŝ���i
6��'�����4�X2#PDXҭ�/�,%�?��� +�ii0�P�21$z��]hک�Uq�p�'���j��=�Us6��n�*��ؒ��M�'9F#J�����Ѝ��J�Wҍ��˵1S։���<5ÁwQEߩhe?ug��]��2�;t㣚����گB��G���)/e���5���{�^�a`ee��P����DBzڧ9��q�F#�6�g���o��g,Q�`u�])�X�m9�v��S�<����߈R���캢�rf_�o��� THז���'ſ�$J~g��:F}����@g��3���ݑ��}�1�ӟfߦ���6�ϟ�f\l!�m2���8�W�0��&^����v3��������*�{v�-ǔ�[���� �����\�P�����h�iv��6���%=�y컲_=���ﰆe.qe�=�Z֘a�6a������h|��y �~��}�6��W���(����$���C�2Q��_8]����rݏ��Ò�1���?�b�I.)��	�@�&�'�T8���?۸�nΞ�Kg3
Q�u"�
u}C��Ga�� 5��/����]ƪ#���ܛ`����,�l�5����[w}�V�ȃ�A��8���9$8(xh�`��2��T=�_��q�}.��i;�.Y"۬%Jt��Q|�"�*������ҥ.�u��`9���-�֚��,3b�)�ڦdw	��4��l�G'lI�@?}ccH��
W���5?b���������Y!�c*`��0��v�L�; �)��F��:�ˮI��	��eF+���	B�nH׋�!br�~V�V�8TƳ��T�J귿�g='{ǧ#���m��	bZ�n���(-��8�x����|�7:������ۺ�� :O>G1ZלuNl���+>������H��^�:�]~��G��Y� &TW�?PF���	>"��`�8��0�y�<�E�J�#��_4��8Jm���w��%��E�d�S���ڏܖ�B[��z����"?�QxE7)8kno}��l��9���*#d �wg�q�,�C�Lx�����1��-��6�xˡ	�g�M�]�g��t�9fG�=��g���M��RxD	�I�]8"v���+>��9|��V��5�g�R�
g���}�;�Yj�d�'��
(��j��oW�.9�?:p�Z�<��s=�^����{n��H��ʔpY�p;�Y7���+�� �b٤����,ˉ��tk���gF3��O�'�{�gܟ���oefE�2�s&���~ȫ^*�nw
����&�d����2#Uʞ�QǓ�E6�^�h|���tbq��*󿣀�iXr�J�0k���z?�ը�z;���f�w�F�X�JmC�tj�?�zC�'_�z�X��myzc�����-��:����Mx\��PG|��Zx�U�rzXpBJo���Hh[
���;���4J�7���q�b-Ta��&k��o+O��CRh�~�h�߉��w�A7c�"Ѱ�ϡY�;�����
��9�}{�N���y��/5��
\��4��P��Pvٞ�͓�A�jL�,��p�T��l��E�Y�%�xh#W{ưԇ�&��O��b�h'{�}��)]�&[�:��^��tV^�H^���R���%NI�R��2P��:��)�P��#����6Vh�/O�s)��-Y~���N"ZO�FY�뇄%��V�UN�{Uv�����`=/*`��27 �����9��t����g�kMJA�)��oH�V:�����'�؋�@��+"�����Y�ހKSd|O��A�@bh�&��o��y�՚�cC��tu������F��A}�%�/����i��l�r�����~�u�O��.�c�@ �#	/i�B���Rw&r�#���ze��má7S����z��uC�l��r�HY�����E��E�Nh���i~0o
)Ya��A6o/��`�/sT�E�PT�1�n# T������A=p,s���ٿX8�(Ow-��O,�Anܔ?tV��ͱ���������Fw�vHr�p��i\N���VF�L��ȟ=6'OylR�F>&OǗ-��?1�����~��K]r\�~U�.�3I�K��c��8�,ecHv�P�IO9B1wV��u��Sc�������M^uL�'��
8#vs����l���B�BL{���3���dXkw�P֕D�FH��V>�<�a�W�6�JU�3����QvC��'3�'�������}Nl�U��Ĥ����w)�q�.[�~�i�[�#1WIW�
+����l�P�ZÌP������#�0̈�2R9�H@�jztU��?b���r�M�XkiN㏲�Si�)�ŰL�6"����(SɇQ������o4��XS�$��#h��C@veXdL��nKؙ�"��Æ�2��w��njN���O �r$u�I'��h(w�ЈFЛ��Z�~s�~��ǥ�ˤ��BN� ��&�+�.%���z_ޣ�,Eϔ KG���Y�Y�$�����(�U�NJ9�m*V�}o��Q�,������T˞z�i"�J�7E ҭ��E���J~ܣ#ݢ��m���L�PW
z|��е�~��Ɏ��='�U&��l�y
�9�k�zh&7��ph�2}cC������ѕ��T�t �	܋�Ġ��ۼ�1��Gtq�<
�2#�anϰ��a��I���w7��.���:]��L����/!:a��$���}#�FF��
׬�0�L��s\i�����p�A�y���=��M���C�<���_��<�T�g�s<�ix��^3���8�.�{̸C�K�E���PVaB�y�@Y�/�+u�U���?��K=����u?��5���M���7�&��3�jd��D�Bc$��4�3�	��Ϋ����ӿ�$Y�ۗۖ��+f�W���y�������Z�s\o*-!�\�-�>��X�t���e���RU��~�f���������e*�P���DPq��x��.����Ϭ|�-����F�6��(��W��=���9���{b��˷G��*����:���N��^rkS��V�� ��Vݕ�Q"�ee�qGԄ�,��B�=s������8뼈'��7H�,�.8��" ׊��h�fL�x�2<#�����5��һ÷E�f��?�� q�|.�����m{ wƭ�l�Pk������I��S�R���A��-]�Y\j=���R�c�CQU0&��_��#m����,o��Ck�ث����=��e����_�`ӎnX�{�t�ROœg�	}������o�!F�t^ �As��R�{��Kt��7y{~�Mrw�L�;�G=ʶ��Æk�j�����Yn�:x�3p�a�'<�u1����B밪M=\<o���
��V�)�|9�a1��~�?_�c>DP��v��zr�����r�؂X$ʅN�H����׃�kj@Lu#\�Y:K4w��_	�4�axy�$-�'BiJ�-%3fir0`�4/
���B�ؙ�,���Q_��'ł��0������A�d���y�d���|�봫]d���plXwF}D[���O�:uP�a�bc`�f�ȼ������G�j]����)ؓ��}�!�}���r+�Z�5�ž��r	r��8Г>��N]=k���]���?!>���&zU�	˲hX<��\t�U�F�	:v[����� I�1�9���}L��5V�Ѭ��Ղ�1Kl���s�y폇:c]C�������u頫��&�1q�/�\F�K�����Q��c��tw����ݚ�cJtI�<��v��K�,�8r떭��S-��t����V��ڝ9^�\�Y
>2��m6�*U(�"	���B�vF�R
�'�������Ą�d�5z�R�q���fA�<J�bҖ[���m��@�3Sy
{��S߿��7^�pIN�ر�,�n��{��H/6���	�3�^�w!��֞�+�A?�j �E:�$8�'�����Lae$ct����C�}�����&�����ƝQ
u��d
nqrl�����=�7�v�㖕b2��#,�{2���ܞ��m|��.
�-oD9��y~�ü��]E�d��"2vB��h����>�۾���+D��~S����x�����.ڈM=-r�(�f�Z�^��|���<]S��Ų��fGq�Vf@Hһ�	�����9�&,j��!��N���'������mH�{a�Z��?��I)6k4���ds��9�9�+vc H�]�\��YV�Y��ހf��K15�st����!I(��%j�#��1��[i<] [v�3'|l*�d���:��)ی`�4��m�۰��v��gl!��D��ƒFz3'A�_�� �WO�QWІ�(鍚,s	��Z��W,�R�Y�m�|ftJw���,���Hr��Lܤ�T���biHi��k �5oO&k��nyh�$�����54s��s稹u�' n�`��'�ݥ��K؂@k�ϐ�.$���2�`h�q�ޗk�� �
�]�N���B��Ɛ��Xѯx�����=�����K��+Zq�ʘQ���#�iĿ����.e�ړ��Z�b*m̍�{�wk��94\��Wn�zo4b0�e�l��$,��%��t�J�������:n�^��}�<q����%դ ��]�7#��f�iI��U-m��̄Q�h{��G[+A!���7�/�It��l:����\��^3��@ek�cB�&���f�0n��Ɂ)�jV��<Ԯ(����p/��8��Gt]$�3IrdS�̣u>�u�?���j�/���J2�&���}ʠ|�8��-�S�V��^�fe�*���������f8K-�4� ,c�Ѓ��k��.�\T��ؠ�a����
�l��PC�_�'ظ�`�-ue��_`.�O���aǱ�]6��L���ݏ��Nsa��+�:K`tW-��%{jy�U�LsE��P'm�K	�G�De��@T��v����a�~E�,x��m��3�Ӊ���9��-�q�wY�1���73�\?��O�0IS*���O���L��v�S�� �aC����5�7#��%��&d'K����x�n�|e�JUd�~���[�����M�U�Wj�zcd۝�:^�(_��r�9��c�N�Q/���!��=��_�x�ٞ�R��µʧD0%M�_"�>�Y{� �9/�Z��G̋����H��z��ٌ]he`q�8R ��⩒�N�-��|_�� wP&��jeG�GK��r,�Bi쑁��R���Ǣ5;��2յ#���?-�@�A뷁b]����P�M�� �j��q��rퟔ9B�8��S��rT�F�[ ����W��m��}�M�!�.��vk�a���'tQg�#�y 8��<��`���#���J����:�5{M�Gl��I�hDObH�	��_��$�����{�[�u���;z�r(����'Ġ+�RA�1޳2Q9=
Cc�J���9NM�Kgv]��k/��l͍GB�����X���5>��S���1��w�\x�/#i�q�D[Γ]X�|/l�搜�KR�����9�3c�<�o*E]��_��Ye��p�\��P�Bnΐ-��qO��@[��ݖ�C=w�[���jk9����c�5�i���2q�Ӯ�}��V �_��lX�7f?`��K���U����^�ھrǟ���B-�uF�`qR��tTX�yD�ê��	 ��W�货�xkI���(�K��䝷cAR��wLyC&��8>���s�h,�՘\�H��ŝGk 9�,�9�`+o��Ɩ�2]�1��#�w��
�ZG�].-��Zʑ�|q3*�\(;�D���&�\�@�@�b��H��$����lve�Q�|�C2W��:���"�"2�-�[�M���#��t{D�$6$M�"������ba���Ͳ���og���L�0�S���Ժ�o�8�,��/��&��t(���D����/|.W�j7���qM�U4�&�`)�����V�P�:���Fܟ�fm�I�e��V�=�ũ�!Q%Bd�7X�[f��2��u�������K����/J�n�a�	ƽ��*���w���Xɷe�������6^tHG=��ƶ��ȷ�?�Y��3��W$���%�2Ґ:���Xp�b��e��8����8���ӛaW�Y�Jn�2�?��T/�a��5�ex'�4FN�;�si�t\�V��Ar@ƚ<��Cy��.R�z&SGJ�b���}k�H�����ق�	p?g�Y�W��SWl��%Pg>f����@�C��z/S�)����Ht��Ġ�'|�(�X<��yZ�
�(��_ڕ�`��R���	�v;"������t��l��C`/�����0��Ɵyz�����q���b���!p~c�Ǘ�� �g����!���z�#
i&tZ��A����zƙ4�G��6�	�0�:d�	�68�Ms7lipJ�RX��$1D7�,��z����������t���m�=�~�� xm軴�߳�ޕ�S1�GJO�Y~fNw�?W;)ʶ$G9*���`�X�`�z��{9_�<�����B��s�/n��{����&���h��>h_�^=]sU�L�#k�B�m�,�����P���y!������= v��޼i���v�Ѭ�c��mL�u�/ߗ� �]l���Uvg���uB���]`K�~JTg�0���R�ౝ�Z3QrK0�3$+��-H3#z�>"0�$�$�q�V?��5u�������Sց��`�<08�ʆm-L�V���Gؕ�vt��j�7E��bw�aI![nw&@�6�~��[���ۇ�N|�-2����Fz����W�L��$��Ӗ�z�Ii���%�^�Q5`{o~W�v��d������q`��L���x?��(�{�Mm�q����o�����ϵ|7�:^0��e��N�PQb�=������ �3:q@�v��l��C�@C:�Y���	Ä�A�@��� �}�!���{U��L�x3��+�t8��wh�Z�����2v�'�0-��ع�]��N�	���G!��p�v���pK� ����ޙ��  {E[���	êI�e�Or���5�Jp�_���g��6G4�pz�Ğ~�z8��K����،}��2u��T�t�E�������1G�կ�J�$G�����.Ln�s�l�����#�����߸��䵭1yqXg$��ƍ��v��{�着��O�w���m�~�<$IW� �������G�.�xO�5�$(���R��^�&������c&4I��AQKS"�=ܜ��	|����K���xɯ��T�$�I$�L�4��'hfCy���qr7J`n�h6֏F9�b�]��"�6��?��9Ml�	��U�p����x�6n��j��1��.�Xڅ�)��N�L�	?�2���*��x�|�H��/0�p��m3,ź��U*׈6��=��#�f��Z�&*�=����o��ײ���ޙ�3����,ǬVW%�> 	��.��4�,���B/�շ����2��ѓ ױ����ZJၤ3�d�� �p�Wo�!���Ձs7��b+:F�mr�f)`�ֲ2;0�����6�Q��	�[��0�'ׄ�=�o�5��M�H��EbsN��tL�~}9#"p�¥���r�Bh)Lx]�+�j��LJ��#!��E(�-�a@$���� Ee�����.(H�RfL;���;5]�"�K��(�fU�����%r��%�"W� ղ��y	��RF���,���h�km8�Pۼl�MU��o�R�2�7�I �����r���������dd'w,� -�C{�����n�]N#Dj�2�>l:��F���g��-`�E�x�<E�$��^hL��RM�p��w�T
�W��$"�;���!��wZ�m�ߓ��3�`�?�,ɊP�n�*���!,�'�:�^\vbJ)�B]e���L�#�����JB����U�!~��Ϲ�o��c�
�qO���Xੇ�6smէL�g�r��k��B�|��[g�I3Qk(tJ��-i����ͯ��~MRT���Q}�N���<�	0//d3��"��c�r���@� �{}�L�q�]�R�Nþ����/��3��j���<�#ru�E\��T�;�o���L�,����u� �&�+E%��	��QL׍�����C/K�t�[��O5u���$*\cc��,MK���D8_���jL��d�O�'��0-<�#�1�
8Z��i7�PE����k�_�(�+==���J݃���.�
�[&Bϔ�⼩�R�� 
�<�FO���d6���N�c4{s�Czj�}��eO3��P�����l~�P���:��m_��Y����]:�M@_���p�m�rx��N�`*]	C��b���{n��Ӄ]�G��wC��t	����fq0Q6�@-�����B��3d� r`���/>A�U5�Gz7���)dā����~6گ&�J*�Y7��<��0|��>f�R��u*M�mR�Ɩ�`�x�I����[���Q\H}���;͎޵�\��d7����%��*���֩yw�{ڌk%P���@Ln@a_��#h���(�����)�}>h��c��[�iwx����U�IJ�lb"s5�ge�m-)�%��R�r����h��_��&ǄSp��y���>Y[��]��*3[�V��b�h�F�.0�9] �Җ��%�4����C��l�T�'�y7�L�𴙳 <_�@܎�\�+K���K��[�/�}��|�G*즟�>N���'��TQ��@?#��Z|����0{ǵ���}8M|�P��ޯ�8X^��G'�]}�n�����H��X�F�uJ��F��y�!�����:W��}����Uk>�3��C�Z�H@��)%S
w����́?%2�X��X������	�]�p��}QUE��v�`2���d�u��I䱳$�rrS��Ǹ<��`���2�gn��E�M\�L�5kT�e��B<,�͵$(�����o�n��[��O��Y#o��%+U	� ̢k�´��[7�$�1���Nq���c[f�֜��4U��rC��v�P�XH��Λ.,�������hDO_�.���A)��/�� �r��k6�Q��,ї�|�ML�����)$�p�=FhP��n,��RC�e%YN�J�<�ٽ3Q�a����[���v��� X�x����Z���;-
���#���.Yy��o��R��]H&3�v��|�����K6��6�G.)%4d��O\�S���(�Y�p����&�eJe�.EJ��x��w�w�l�X�Pq�y�*@;�(4���:��;��v�9���d�C�G�d�֏����Q��8��u�@���w\`�bc��1�z�~�H���0Ą�p��b��z�:G�s�!9���>Wꁍ&Ju����pԫ ��e8v$����݈Q\G�����s_�5��N$���w��k;�rR�ۚ��$��@	o��o���������
�y�R:�&��"/�E� (��4n�P��cs����9�i\c��1�8�����f�R 8���7�~'+)U�f�,<����;}�U�����UAyL���1B�F���oR�.S.�c�<8y�znϢB�q
.z���{�U��^L�W V�)$�dY4+3���8�1.&�>������1��'>�?J�y�+��O~�;�ÐAR�����%�H`zp�{� ��y�1]�c!�sޫ T�&L��Ǖv�/��*��2O������L��tx�ܑp�4�^p|�їuЃ�L���HWQ��D�*�`�%�~��%>q�=�<$ʴ�5��i�yj˺hEZz��w���l�9�bS�V����'	�1���^2n�6e2up3�X�q
�޼:K�ҷ`�h�=�!�b���h����:�u�C}sZ�^���w���L�v����Ƽ�&q��_[�t���h����P`U3֣S���kB��o��f6'��+���oe]��S-��E���`��?{7�\U�z%@�!&� �����m�=��&{�,;���2ّS�]�D���֮mRw�-�������TKڊ?�
�׵���*���y.ș�-R%"�t���Z����o�2oa��A��ݕ�
�
q�4�J;Q��ዋIB��3B:�f3i��s�!>5v�a�']E�Q����6��np����#K>�4��}4 �E-�
�C|,��^L�<��
9�"������o3."�r�4ҙ�7(/�9��t���8�5��%�X ���|��W��WL����
�K���(�F��g�U�ƽ�v�H��W�q�a$����%_���᳾���'��Mw�vyλ�LA��G���*�F�8{m�F�7�v�W^Ư�jo�g�ʝ]�� pF@��"����Y�D�N� �� 5���xwQ@AY@Z����1^W@�.�6c1��j�o2�P8�L�G ��G��#�iq{��I[D/��]�D�W+�&#����lhbe�D*Ɯ[�kJߪ��c�}�z ��^ �_�~�xQ�n>��&��)�^�jQ���d�*�����J�G!�)�Md����:�����Y�(bd	��/��I^o�4�¤�4��G�N[�ΐ���{k�a�f1�o�I�EV݋1�W,jS��%�;��n_�Di�8�g��{�~�bC�3V���`t�.�ս��t����2I��e�����6�_���l \����� ��:���WF�z�w�pl���x�4	Iީ�f�ĳY쯂��]������i�m��@��W����/��;bx��p�i��1$)�8�&�[?d��g2�'����.�ѯ��:����X>@B ��V�K�o��'�����4sߖ"�C�E� *�f]!�x.;���N��M��U�Gᔨo^���;5�dʸ��G ���Н�kV�ok2_z(������`�a�a"j��N��Z���.�Z�,+�JW/�"�a<I'�a�T1�V�jz](��ߨS�1>)���^��vF�j:_p�D��m����b���5bc�`w�:��&<�����<��*������gb��Eŵԉ�G*��
�[�Z�R-"�M)�k�YEKi�$Z��y���ϵS?��z�UB�h� ��9�YL���}Oj�E+�t�[��c��J[O"���$e�i�ʽ.7���	h�QuJ�F�����TVut��)�n�%q�LcK �2�;��,'�h����?��L����l�sl�Q���>���$�K��m(���Zϓ�}�MNFM�Īy,�g���aIqB��鄼�ݼ�Ц��f�����*�Ǒ�K�c9G94��>|�q�{��e+�MAЭ���� :����k/F8��Q6.Q%�T�`9>�r䁺2ԗ[�tO�V!�]z�:�U�[�P��xΉ�r�c&hQ��pn�F������46F�ZY�̳L��4ve��65�ZȌ���y+�QS�����T�L�#��8�`�F�nMw�~`5��a���B�C�<�_�@8��g �
Yt��w�?B�q��1���lJ�s������ɩ.�[kL�D��%����& y}�l�P�&�y@x�����:"q~�t�O��O�s��G���ҥyK� � .����p���06H7�T�S�]�\�U�P��V�*��R��lQt�1��=��P(�+��n�E:�J^�}Tt^'K�ꨒ��[�z7����	�H5�&���t%0i�r\qw����{�Ojr���/���([#�w�Hꨂ����rXg�9�H�x�΁sL/�c��}q=����X54�F6�&i�a�\u����Lԃ[ř���G����|�&���_�4�%#�*n� ۼ�΅p3��mcԾ�n�~)�8��/cT�����n� �US'�A*;*�V���-!�Ӑ����@�uy�� [z}�Ԧ��mb�(]9Z0G���7��)'�-�UB�}o��P#z�ʑ�Wě��i�
��@{e| N�+�\���4#������\+ҦT+�'#�r�%�K��[ESfxŎK��z�wg���v��W�11\?<�Vx��!~6Hڶ����|O����h3�Mb����͌�Pc�چ`{$ɨ��B���J��Kz�ND���HɰM����߬4�� {��A�'�<r�z�����O��3j�} <ʲ�B�z�N�ꚡ�2�p^�0/py_����u�j�� �]�(J�&�kiJ|�������iBN(��`�W�1��6}�j�ô=x2�]�'T��ֽK���0hC|�&'#��7{�	���J�ϧ葵I}��I0Cz	���ua��@�`l1]�y0����������ܵ��R
��	
��9�E��CM�I�6d߽@�'[ɱH�[f�d= 9 �9��۲V&E��~X=L�jyZ1?):�!7q�l�ٕ���V����`���^�dbI%`�ZH���F�y��6�k�g=�}L�]�ΠZi�=���|��.���8�4�O�5N�ٹ!o�c���3����7�����SG�jf�����k)(<r�L^57z�^��C�"�Qo���\��q�(�ܗ@3��%W4�:z�n�FmFM�����6���b��%����+0	Y-¤@4L���d��������٦"��su:K��6:q��&�y랔�E`�m"��X��#O�h#H4X��n_�4Mdzv����k��EIHڴ�!�_SB��/����Fw:/)T�J�]���٬�+�������������ԩoc[���=���_���ˮZ��x�m���~���$�k+;h�O�L6L��e�u���k�g����1^7�Ʒ�b��2�s!�O,�n00}g��%�˹�5V������n�/���y�ޕ?9G�[�ӻ�m/���:ڢ��[}����qΦY��t����gv�y)��@b��W�7��T�#>�ܴ-��F2Km�51t�0�`�M2��8�Y&�|�dR���7�C�x��CW�.Fc���y�Q�+.�����{vO4�X�D�s=M�|�	$��)�evR���zu�jҨ�'�(�����3=���5�㊓%��=Y\ԭ}���g
�e5�^��F$�;��ۡ�X"�l�bL�Po mR�0����#�pz��
��q��0f-:v�����E�ǖnH!�0K�����6F�
��7�w�� L4�J1*��\N��BPwʡt��\Z�(o�}���Q�0΢4Wn���Bb�1K����ׄ{W��5|a0m'3��x1}��0��N���0��~�ϑ�Gxjۏ`=�����o���_׷�d�`g:-����E� �w�Z��=�L�� ���z�@�ߢ;��7'��h���5 ���̸b�$�<Xig征�z����х0��\_�AW]�u����W��;؝��jKuh
�J��|EN���,:��Y<"j�?�<`뉘P ��Q=�9���P�� ,�y�)̪c~F�ݚ�P�z���sa{u��\�L&�z=�7K��̕����o������..��^R�y^Q�,�tlM�s�u�U��ˆCe~Ҧ3�(�R�(Qz��e`�U����0p7���ML�̞	2P��(�[.���s�	�W�f��T���̐WQ�:o�����xd�ڛl�e�[������M�m��+�R-M�b��������vsvuhUP�@Jh{m��<�vH�+WH>��I���:���W[�x�#m+B�����D�ϗl��ljY�Nu��rX��J�L��x�k���Rel�W��N@���MvE-~S50}Cx�����ʶ�u�Ȟ`_G�l[�?���t���#tj@;��	�T�V+K���*�Z����5?��G�U!��h���j��x��Zd�%��U�A����l�6�N��br�Ѿ�r	iD��2] �����5�e���/���׭��_QG*�]q9�k�Z�T��kfQ�'��1�f�"J�J���A�D���r�g��!��lZ[��6[9O�a�;�_������e�E�>���$~��dœړ�v�@��Y`l������1����E����| h<�m��D��
�Ą��h ����/2�I���
�}KK�`r*?{��~
n�I[��}�*H� �uadi��ï8�n+϶@�"-��c��O�Z���b�}�Ճ���Z�s���Վ*�=�Q���)�8��,�?�;��>�3����B��w��T�AE�S�<�M�w�	����9�*��u�B�6.�Ɂ|�����!6}���"�ʧ�_U���nI�������_�&��+�������,��OY��ܞm�{�9W�u���u�p�-�7�Ew�JА�'$����+t���Uu��]�<8�����f2T�?9�̴>�w6m�ݟMG�Zu�p���dCF���� ��D�Y֚�ˣ��i]%�X؞�OYHd�z}�Ǹ�����+��ʠ��|jb���u|����5]:g!���(ss�� ��Ϥts��a����b�=��3�v�#C�Z��T�~q�A��DiѢ�dՀ�����z������/Z�eO�Q�n�0���֜�iLb�9Fo����$`���A<�ir��qP|���������`�1c�L&�6����\��ׇ�jV*�IoI�t�G�����u�y�z�H#��?+�
C���k�ڃx!�
9Cx��WN�z:�����U;u�]�A@׍�&�R��b�х�܈u��Ї���]�Lb|�I0]���3�;K��T>I�YaCB��s�������ʈ����}h��9�iDu��T�&�Ȯ�VV=h����=R8��)q�V�d��|GAV1NXU���v��3^m^9P`P�8J�������2b��=6���4���sWyᏪd��I{����&p�E"誴Ɗgr����t����)�2ÑZ}�����.���'2e^���M�$��.�=9�iU�K����s�'�20G �
��-���������[�����0o��b�R(��S
��_�54��E��Cq�ɜ4�6[O�/U���c嗄p{�������2�u)�����iď�"֐���	�_lL�R,�!�(��!�����۸������V8�q
�$�r�䀚(�0c_SH2���u�_�ܲM�sDǝ�� U���t�=-��-kٜ��a��@�e+����B����v�����t�4CI*�g/�\� �"Z�=��B|�m�L���Q���vp�!���|�Gj�x0"�Lq�>�y	�ú�������Ԫ�M� =��eʁh*�B5͙����'a��H�ʞ�`�_�^q��S���l�ePV�/ ��/�K־)���B��X�C�q�o�q�1���Q�З֌�_��.��6N2b@n_����t�__�u0D��o�<���!�^���nLQ�ď�x|3������3A��X�<����*�F`>.,�u�3�ClM����Hk�}*Ī�3XnV�cx��@~�� ��=�}�	��߄ k�o3v�u�|�"ic�O�%�B�R��=���xI��M�0�ғ�6~v�@�AB1Z��+v�;m��Si��8���F,i[f�6ѼD��ō�K!J��e%to7�0x�o�y���.�b<O�%O�����%5P�p��?��y���?L���ȲŰOH���D��QYW�{W�����^��B�������j�U ����ش�;�o^�V.���t
�7�|^��*����NH��/O��cxM@;���T�!�0� |����B=�*��-����3jg�����l����f�����M4��O܈l.��`/5@/�9�+ߖN���6���;t�Ϙ=4��F>x5j>c�
�&���4��"���������>�>'4�_���X	S����Hײ�'m�t�̼a�1��v��h��^��6{�ŔƾMi��5͵	p���"M�Վ��5�P�鵒!
�?!��Km���7 `����æ���|�f����~��m�D�����&-O�B��
�.���;��X�4�n����T���i��Y��Kµ��`@�~����w��d���e�RVr[I�P��v�aɠQ׊&��C�gә�P����¢59�A����q�:�T���������u�D0ىK���Z�V ��8�Iq�R:�ט�3N_�~�)��w��l0�Ć��ݭX�������|H2�,L�O��e�R�C㸪�'�-\Ɂ�Fc�4?�s%;��D�1|0B��TC��en�L�i��ת%9���hC���J�4 ���[.�ҨYC	^ۨ,�L����\i
��45����_�I��1й,�����I_1OԲ<-�d�U7�X�'R{�����F,��͟��#��_���i�4���83RZJ�Xk�� ��GT�!S��s��1�x�v�~��*h����`�C�2�K�Jx$��kKɒ�6���m]�=���M�M��^kN��[���0�4�c�csnYb��)�d��⣲AK�"K�`|�L���,���0��X��EO=/�p�{5����>ÆgS��� �[��j�wKV�!�zQ�  .M��Hޤ#���q��3�γ�MV�������8;�,�
$^�H�!N)�u���G.���EH2ݩ��%��s�$ǝ��
S���/�^w����t>:W��v$�&����{	{_R��)s�F�2O��J�~�\�j'W"�r�A_�o�빀�K�>[	� �ci>�Ĝ��f������sV�����&�I���N��x��-�\�GZ��=��L�
/��0�V�}3O�n��e�VIv)a5M�$����wR	;�&sI�P6�]`�eOHN�S��+�8o���x;7�OI�`�D�R�d���Zy<[u����cBۜ��]��@�Pܯ�KS?(�iJ G��k;�И~�g�E�����.��'o������-�/�;��[�[����9����֏���W���X��*��$�0�E�X���D�^�r{�D/�ُ{��S'���X�K���V}V>n5�P�F��uxb�8) z�0��餍$|��L~�0�!/����Z�9K��(ƀ�Q8�n��F&D����n���T��>�4�Ӡ��Ĉ5�]|E��k����2侎*F�����u��Ė�����sD��A�a,��l<��/��i{5��ސ�}�ᢂ��_6+<T1��"I���\�Wh���J��m�m����r���!hh���'լl	�R�#ۤ�#�@\�B-� O1�U�
pHI�OX���50�K����&dga���>@�9܌��8X�f�N"�]~g����"c��q�`{�K� �P�M�e�OWi~�N��/�Y�X	�a�YX�ũY�)�+=т=��*]��w����2�^1�5���Bs4���w��/܋"�;	��&��!'b�*����TҾ���6�%��E�}Z��c��
�L9qF-SK�	�s�^��]����Q�9�?r$��C���n�&�����н�+Ѽ?x��8�+���\�	T�r�e����X^��d�y�'#�:�o�X25��\�ˣ��_��Zc����xl�P�K:��4�>G\�>:������dX��8i�؎m���#�\��G%J�]T���eZ���h'.�._Z0ܒg>U 힁e�%ZV��H�MGp8!�p���7DA�p+�D���;�r�*����V�e��t��[L]c����m[ ����Zr������;ˊ$�;��LS��]L{�Ц���̘����6k�����є�Kδ�f���S��*�"�t(|gs��`8=0�U����Ӄ���R��\g.�G��5��bl.�g�V1�{�~|+
��g�spZ�� ��`3ǣj��W�jǠ���@��%�͕��/�.��(��_��Nh����`3|��7��Dk�d�:�ǐ��D��[���y�C)k��x����( 
��B�_����:D�[.n��鐙Q���Rn:OC7�Aoh`�5�GTś�NETQHv&�����Q#�\e�2*[W��v�U��� �W�+ӣ�8���]tD�B1�j��W�p�]jO�y�k!|TS*kxn���X�XX�Z�/dH:�?�v��}�O�-���L ~�)�m$>�Z�[>�k|*4���w1j��u��0�s��!�ռ��j�j'k5@�$�"A�	��:��v�C�,mU@�xS�HY�C?~@��Y���Ge����j"��B�=�|���Quɥ��x|�r ��[9#z�}��8�'�L(~�P5g�V6��x��,�C�?�˘�ʞ+�90��\�X����N���\�|��޵d��*,��|�k��T�̯���0JDڅ�	e)�g)~"��U�4qg��0i�W�G�Q�(���$�I�4J���������VG=+��z���T�'>}�-΀3��eX8���=���{�����>����4�|f���rs�`�ߺ��7�f�I��nL����-Y��U+riپuR�<v&�3�z�矟v7�A,��L��ƞ�{F׈DUIv�MB�����(��;;��}��v��ze�9m$"x&�g��ׁ��Z�GO^�����ԛ�Py��([3O�8�$�}	���Su$�sg2�)�=1�|��5��9�B�2�M�Ƴ{�kg����=m;�8�J�~�(�G"������oJ�[�^�?a�2T��"]Fxi�h�XZ�� ���:��~��n��ŝ�W*�f�8��N>3Z[���sd(����У��*~'vݦv�C6!!�֫��KII����1�@�f��F%NV/xC�K���X�*�h�G�x�	��d���6�ᓐs�G9kd�Ը�b
�)���V�D5Rn��s��>�Mq߀�r�cKOt�C��b"ş�)'���v����+�j�9���}`Aq�;��;��g9<���G����ߗ��m�ϙKA4r���}M�VhӮ�g�r�j@dRc��6=?Ϗ��B�����{��7�Q�	)�N�bD���w�*I�^��AdKu:�q6w�q�N�q[��Ew�꫇*���[U���8��L ���	��>�,b<`:q4H�zL����F�q?�+@��0�B�G����0U1Q4��l��n	]�uղ",��l�-�Z��/+�!ω�� Ex�H"�YD��o���}�)��3KL*��^9����]5����}�\Q:�ݨ��~S,	i�8�5��]�G����Q�X�A�ðð0�" S�<�cY�E�h�,t�w�=�����br��Z]��9D�`���4M=e��;��AdP�j�S/�ǧ?�}j(��D}�8��K�L��� dp'�ל�C�>���r[&PL����0��mHD�;�0��IY�ٕ+ٛ9Ijp����d���tZu���X~@e&�O��-4�մ/�L��ld�Ų;�[��<��S�R� ,�wZ�{<XO��P�gĕQ�~sjJ�<t�z/���)��/Ak��9��v�ך�Dw����h�_Gn�wq����A�N�.�>�
�&���>��ڕM��,�6����[s����q��K�paz�!�"��܌OcM�t��?����y�Ԋ�G��_Vf������)QW�#��HZKR�Gl�G�YL��5�-�tm�{��:��本��h��ʽ	FF�����0قé(��:MU�}��ta���znͮ�����G�3yi,G�J(#��Q:�aD����i�Q;���.{h�
Q.��٨DdBJ�����$i&��������u�z�wC�S{*������$v��`��K��c�&�sf��\;5t��_̞�x_#�@n%���N�Lm��R圾%!��V�&�م~��Q-�9>�l���}&���Qe�+��?4��^Q��biK�O0N�|��� @=��' *f��q�I������֣vtx�}₎Y-�0I�D�Ï7=P�� c�|������!�R��w�s��c,1��L�Y�t����M��.�8ң��o���U��j��#0�K<�K܋��˵�-A�(�a��H��wKTQ��y^�I�4hiD`\�6��1��ghR�^_(F�G�5���)�\���8!
���i�z�{�</�S��6���'J�m�?S���X�w��*�ٜr^��c
��	�z81%�`�ޯ_���KH]8/�N��a����kV�X��틦�����FN/�r�/4�)$OVK?���S�%(hL)�3���
���5�BZ������῵!]�g�:S�j"6������gp�D�rB����x���Y��y�5�@;���`�h�?��E��l�(vX3�2R�û�E ��=ҹ��������n��dsWn�X����[t;a��S���!�D^lY��;`qq���!t���u3`�Ԯ���-�5u�2�mT�U�e#ӻ.�O=�ؔ�$�ơ)+��n�tC.��� y1�^mA��-|/'KXTW���߬"��<���M���l�(�h1t�E�?��p�������d/$[�����\b���T�Y���	=��}�k�����߹λ/�C� �[�dt���#�]�N`��B �X�B���r��(g�KQ�Jns�*���{��mnxơxa����eI���r��M煮M��PLL�t��e,g�b�j!�G-��b�3�����݉���WW�#A��F�$_g�mO�+��t�c�@ʗS)�<�~�TqKxk�?ܛ���i�ʔ8�OJE�X�~SP%�e������X/��%<�
	c�Ɨ���|h(�ښh}^>2��2(���4R��k"}��a-��ð���W��M�Q���	�Tpvk�ԌXi�[2
�s����m&< '�C��y� ���&��Н���U�\s64@ݰ�K�&�l"�	�78qzI��Ѩ+[�D=� b��eVf��˳40"�Q��t�7�,�eBD��9b�g�J@��:g�#Z����"u�Ys���x�נ�X[�UNXй�n���v�u��&��ga�T�u�vi�U��SݕU��=��3Qx�MLU3�7����F�mZ'�	��:�1'��8S��o�kN�C�_*A(��4[��PǽWD�;U���w��cٸ�Q�*
 *��xH�F.$�K�$�L�O�A*+!�	�3pB�a|ś�����,㎮w�����s�s���4.�����u��t�y��qzX��\�L�"�X��U|x:@*�LWĪ?�D ��IG�/��*a��[Q�2(@� �!��*�*+��Y�������G�^�� a/�1�FY���?�#���L��A��=-`��B�Vɾ"Ld��p�xz���pk ��H�g�����j��?G��u5B�&�/��43�)�#�6Yu��f��|��Cl��D���@��6�Z4͑�e���}��R� h�r65/�4���{<����F���sx@�:jt�J��z-ѕ��Dg�j���R�.`�u�l��^���s��$7<�T�����̖Ǝb���wtq�x`����b���i�<� P�C�uM1ݶ�ć��=�7=֠�1 (���q�hhz���^�e�4�_�y�*�ύOĄ��H&�^0�j�����R܁�T]>�[zk"�Ulͬ���+������P�OSskR��㏑*�� �"���D���J�q*�#�<�\�,c\��<r�&��S�	�a8U�y����`�9��tt�Ҝ�d�1�(Ekex���iK\�������y��&�>
��$�hw�!������;�<@�kHK
*��t���C�HC��F}�E�����A����ò����3�����o*��Z�C�>����X�ou��|����Bh�)���:s����B��U���\4w��%�p��!������%��S �z�SX�΂��x�AW���O $������`�	�&��vݢQ?+��v���,=�`1H�S�L��~l�hw�h8�Ϛ]rP�C7���&��0�����rN�~_����Q߿ӕ�>:EB/j��y������I����oFұxC��Dh;pfݑF��2��aϕ����h���e�e��r��z�[;䆎>�)�
���.ŏ��T�r�l�y���\G�RH�{wTU-a�y���f��ڶȼ�mt��C� 7u�Ϸ"A��x~�#�rj9���0�Y�j��og��� @�>�ؗj�U�ȲΑ��l� �%Ooa�{�ڿ��! ͩ�#)sZ�)w$�N�Q������~ƴ�:�l.�����Ü+�i$r�gy$���K?�S�*��#f2��s���!�v���6¿�����(m���C�	.V|���?�Ʊ��*l-E9"pT.��	`:vg�"������WZd]��[����IXL��N���8�7���B����+�"4K_'�Ih�՘uj��d�K��[�I�:��S�[&��s<y���JvV5q?		 ��II�������Y�-�Z1��9���������M�O�U�7�_���V{�I)&??���,��wh뼆5������NRᨩw1��B^�n�J	93�h&��|��}�^�d�}mw�Zk>�
 w��s�u~�D��akVO]7Y���+8�w��M77b�U@�cTK���݂��C�8s�a���+�
�Mg,������~r���i}�U'�`�����P�1N��7��n��g2���XV��+
�/�Ӏ�b�g��+�C�otW�.4]�FU��(��M�KQɻ��N3�A`#q�G!�[ó��!raĚ
�`���u�n"$�p�-�D%߉ѱ�s�X�Dl
�Ґ��>���4吤��r�np��W��WTr��WLa�fo�Ԫ�~��6�'���J�`p�z��K1�M:ly�~(Χ�1��]Ŵ EE������/0>�4��ˈ�-�-��f�Dצ�0Z]x���~�̭z�*M����dȀ��ݴq1��!7��eK���F����ɾ���(N
܊%�ǐ>�$qZ1x��+����=Z����o
1A�y[J�q�����2o���?̑>J���}v���
�=����j0#]"Sw��]av�M��~�ng$#�F	'����gVL�$�{��#�Ϟ��L�����������p�{��l��WvŎ.���=/4�'їfo����hFA�٦%���0�B�1r�"pf���8^�ˢ[+jLSM�̈E\ƺ��r�g?o�wl~��I-����EbT�ò�!N�)��ʛ>k�t繃Ћ��l�1{�9���ti�eS͜�JE��Cp�����[C�=���"��/7�!qǮ��o�x������X�:"�Fp٬;j�i|nP�c�p}�55{桑OA�Jİ�	��*�ꖰ�鿆?�\Xt+��Q�t+)Y�P9C�*�S��q._�دY�n��gk�i�!���B�A���`��`��J�ưa��� pF)#o�*_�@+1x.�82A����1��kJ��	fY,���A^3ODy��

�	�WڧE�������P~�>�M,�����I�/�lV�2 �D��X�y���2�R�������,!���%gW�~��s������4 ���_'�c����~�'c;���{��F'��}:�"�80M_�Pb���E���\h�����ChuhK09�.�9�$4O�L؉���j�<�ʣb����FiU{^��z�˘�YG�E^��GlA} &� �@E���|��7��T�q�H�E����i����#o��*nb	�k.3���{�w`���C�i�O����g2L��ݩ�4��Qq�叧6��0�n}Dz�z�܈��V4��p8�f��,�'��^�|b�����Ĩ�@��I��^��3�ssL��,��i��M,°��L�qJ��:���x�?' y7}�n����?�,����^��L�
�)����n�Y��FB���|L��
�vD��?�M>�L]��
TBmʼ��{͒���O9�^������e�Z�);!��ƹ;c����NT���Fˀ&y��wwd�������g�"b(32�@]K)��A�i�Z�
��Éb"zw2�.Ac���jK��Ŗ@s�P������r>�Pұ2T�@�����[iV
��)�M�Ʋ�����2w$D�ӗ�M�-�E��H�z�$4�/�Pk�F�ǘҸ�;Ɨo=:�o������߃�wv4��s�����dLh[��j �{Ls�2^t�4��Z%L2Z����t��{�<T<ŧ@쁇��眏� �i��V=��<R� �31��pi{�*��^�������%g۶su&� H��y��yH7�7<g�VG�s�\��#X�=6��֌ "�$�"5i2c� �^�G��#Ƹ����[SExD,8��ʝ-�'�_�E9�ٔ2����L�ʛO�?�ׂ:��Ӗ�TϗlMIM�f�EN^q!˜�������Z�h�@�-�߬O�Z���^R��
RJ�g4>����r�2k�C}�P�nAA-���\�D��֫��<}<�(Q��I�K%�r
���	�����P��N���4�3U���R�Bʊ�1H-؇3�eo�u�����	��� �/RU��o
F��Ձ*���&��	��[t���94m���� �L��2{i�?O�Q]r���;�oj��Igo�ҵ=z���Oló��X2F��I�'a�OzP7܍܄��s#V���xi/��u�W5�_u�=�-Z�#�&:7PHa '���u �6
}��43���J�C9��������:�!c s�Ė��ZTK�����C�*}yh3�y�2]$j�PY3~!�<ԅ29���-�x O!4�GT\�wrp1��ff|t� /TA�����nط�{����\��q�k��rq�,�������,�bQ�ǘ;Vo<�ж���5��.I�
���g�n#��2��w�!�:����߾/34~�T�=.����9y��o�flcj�i���1*�?��	C	�:�T�3������W�O��v���4�K-7��'��@{�V���c���w����{Lm��:2ƴ�Ē��~%q�9�:�y����s�33� y��x�Mx��P\���0��L�|�u�tg\�:F9�p3Z���CǷvB7��&�J��
�_�N@cjc�%=�����.j��r7G�aO�d���La�L�To��e�N���D��pL�������J��Q��NJ���՝2�K�(	):!���x̘ӊ�gx�����LMQ�E/���$�������I8��O
b��/|�S-/ʝ����	;���hg�߇�섹�y1�/�;�yC�~u��ďY�vv0i�m�Λ#i�?<�4�A������h���Z��r#�����K��H�z"38G�[���@��6� �I��M�q�� ����Qu*z�GzxPAݓv��A�n.�t�4�Rqv:��	?��{Z�\��{��R'_Z���V\��l����6��X#��r3�j����;3�q��Q�V)t%�kߺk�)� �#���W:�v�e+Sj�����,��[&[���n`�]q &HO[�R���z�!w0�Q���n$B=��IƂ�b�J��텭
LoL��?�4�r�����m{�I��k*?�C�������<�48�$%Y)[�19�X#�%[<	�V�&��+}��NY3f�Ok"-�������&� ߫�4�~GF�<+,Zy���V>=oR�#���� �>��q�
ܹa�	�9L��3,n������gb�$���5���J��y�*`��C��m��L�u� �}�"Z�{�:�*�`�7���1���xS�C�L�Q1O���pG,�ˊ�(�*b���-���>�G���7�QH���)FG���G.h��g���L:��Cv��>[�i�r(v��!�Q�7�i�^o8��U�7t7�>4��H'R��(�'�F�\�(�"��ɑ�:#`�	TF��;uX�	�S}�弖��k���N����H-ڠ���J�m ��4˲����c���dy3qIfk���$Z�1�fmꀑ��K�@���4���<��~tӓ\N��O)_��=}�/��2G�t�\��JMg���]��< ���꘯�r���(:��B��.a�j�1�ɑr�KKZ��G� Æ�v��g��y���	�g�p�:���e����yŭ�g��칡��Y�0��]��tB��&����/7�V���gW��p`���GC���A:m3��봊����)�q.d�P�Lծ>��Q6d^l�)��D��Bڎ/��,�Rk�\���e�]�y��a﬌+T9�x��� xbf�0�hy3�������wC�]��[��=���tdcK<n��&F�>����c@�a��x*����H{@��s��c�:���o�
=qZ�y�drס����@fO�H�Dx��2�<�~��cM$��AA��dR��~S_�J	�f^/��y������#�f�D��Gg\�c���Uc�咧�	ۥ�)\_8�\I+�;%�N�!w�	ݹ�5Ю��8)ʓ{>���!ۋI��#k�r��9'�e�������\�P��1&d���͡j�ߙ>�����_��9�u3��0T8V��uYK7�y#��:a���C�Uçd��gPcc�́	I�����:�����I�g}�ow�`��Z��|JP����w�Xƚ浦��䢷�����u;e]߻M?�[��;O�
"���?��̓�Uyf���jϒiL�t��|��y���Q�������!y�OKwn��M ��t��z����&^�_6h]l�6�Iq��S?�T���˃�J�C�p��Y�U s��"�j]�/�z�NSb�C��E��fa��z�O�O�;Uf����F��%1bM�<�1X%d_�S��Ü�6���!S�߮����0ı_Ä�Gf)hMoЁ�ϜF�ͼ�aW�D��.�y\l��H%I�)0�K3�|��_�q�d'�����6v&1��7mR;$9�<��S��|��d-��v�L�ryG�9�éG���̕�٥�/ϑ$zK��Ψ����^S.�>�c3�#xR�;".�Oi������Bώ@���L����$he�.�������
牫�T�m֕��1�EnG ̡���LDPt9W!r����2�3݃�UE��
�����B��w����Ǥ	��}�פ�z���P$3��t�=$�V��kv�����G!��3�\v�@�_�9O�c%� �1�c���ۧ6���0j�4.�;V.�U�DI��}��:��7.!���:�v�����ݮR��&M��+�0�mU�_�އ�,��iX�s)���n&=8��X�HZWؔ��@�9~��)���P�"m��y�E�F��J�ʮS	ڢ<uq��	H/H|
mI�?%:|h��.�K�5i�n�+u�W!�*�L3�����X4^��ʉA4)�ul
�9�#!֌�g��Te�����/�L	l��Y��)e���V�Y��a�����׷���i �vpl�Lu=Ow� T�F�EN[iq��ܚ"y�����V�|�(�}~:�̎��0Cu���2]^2�zԗ��h$�#ΨTϙR4|ϳ`�x��Q����P+���S,�
�@�}��8�$ ��0�����U������$XQ��}��LA}S�B{W3�?A������>9�G����x99��1��'+�6�%�q�%�D9X�/b�\�O^F�)]�`�0gX{�?�+ކ�%"�F�x���}�j6�h�7�1N4ǮH�-~8k��zvb^�)=#��gK�}���ZЀ�~#��J�n�� |{�^צ )�.Z�?s�D���+p�D��7�.�<)���P�Q�3ķ!���|��Q�'t��;~3|�58������iU|��b�C���6{֑EꐗVO���L�yx��}X���-}�֧�����ѹxA��!'��1��^�C^�cCԳ.�r�TQ��<��Q𬍊�j�����%8�}�:����?ߢ���*�t����p'.fr�Pu��MF�,|$W$���"���(�:�6 ���Y�y��!�	���=�����$82߃���*_�	����B�n��ÿ�Ń��r�,~U�O����_!	g9j3�S��2�(�PNfJ?A��1�BhŸ�]	����9�m/߿��3��9�G\������-���tK���%�,P5�h�k�U	Q6<cto��V�j��]E��*���@18<&b:Վ����v.�|��^��!�µ�K�C?m� �Ǣ	�o�|8��L��y_�:�M��R}�'n��#���ư�v`�J$��T�UL2n��$�I�䊠T�� Sg�rr�g��j>Xa�t�.�j~JIcuZO��S�4��I ��K��u��k1�n�%���c%fG�:}ŉ�D�nWZ�%�,`�O�i 	����o�	��'��C�z�S���.�j��1��ڟw�5"�;�X��J}a�3�N�7��f�㿩�4�`���N���zJ�n�h Kɚ0�y�Wi��q���,z�w�~��_lcjHNM+~+�Ѩ�[����Zh ^G��8�F�J&?l*��.�T�׼��L-��c�TCỺ\t��y@����F�����B*�nCh�$�1�''E�'�lͬ�?����
ʄԪ��\�!����9L��j�KHoK���O/4�ċe���ɿ_����+�z�s}��)�MRP��=����ϒ?5j�z
ȟ��B9�8�&�{��V'�k�X�o]�u�}�J$���_��+,��ғ ��8>������lk�p�n��CIʖ��_�E���@5�F��<��)�?Å|������<B�U�R��E����E���%�#����	Ȣ$�*`�T�I��&yG�F|���e�����T��!�u-x/��[�wDI�,�"�D�8� 4os�{ֽ}٥h�c�<�Pt����I+�T<�5a�Q��h�s�K�+�#�2����Vwp�j��ŏ6�!��9sa�����j�u_��nͅ���	���T!`��+��^������gĿN�gz,��b��jkz\@"�P����_��e�RIf���������U�ಸ	�m�[��@����������:Ɠ��s�Jf�F"ռ�6̧�j�Q��`r�n�����:}����@^t�a'�-�7����3�UN��*=&�2\w�f}�"� ȶR�0���92����S �B<\&f$B�M:1l	:�T���2�r<��5�f��r�J6;Z����X���%j��R���n�Y�~�0	�C�0Y��H�4t}��WEe�nF@��ӳ7X�BM	1T)q��x@���g�<T]^�����+R�^|�$"^M�����Y��,�Ww���;_��f�Ud����A{�1a�A��;�"je	�����������A�9+�C{��bbf���'U;���&�أO��$.h)�����S�$�V��"���!��8`ğ�Y[����Y�I/�-o�6�b��h,�~UB��f� y�Zi�7�~ÞYܪe�س��&2`��[��)A�Qc	ң9-�6fư/��̍�bҺ?���Y�Z� d���79�a*��Keb���8���R�)bE���Tw���C��ͣnP���'_��_qb��CK�/�����ʖ�mԏD�5�a�3c,�YJ�V��w��9,P��1�l�t�r�6�AgAη��R��zu��P���H�!'��=�B=�S5IP����
:М�*�0�ypcm�{��l�`�{����I���6����d�1nX�$C��Ӫ�u�I�G"�딌�����@^�j�<sm����c<���x��w�T�#�14-ˋp�ȭ��o.\k�l�/���K��B���]g:K��8��<G�g�����9Xgί�&��	f�n�g�Py3�w�5~��
���U�b"+�xw��^33!a�0Jm���w(
4s�yσ�g���	X�ι���0Q&����¤���\�&�nG�:����p'l~�p�6ĝɢ����;��$D���Z�0ܚ������4����Nla�Uh��#��V8K2p�]n|o���+,�������d)w����b���w�|8��%ڂJ�R�U�X�f����J���[�*�k�m��M/��&u|o>��u0�53E]�p�y@@4+�y���VR��y������:3��fQi��k���-8����]��FF|,�U_Ш�<*��>c,�Y�ƒ��߂P�����Cg���a��I�^_��-��X��T ���<B �,�(�4�)@?�D��wq�q�@�6ݽ��gy�_���d)�g��$w(	��9�]���۶i�=e�<z�7�c�nfb1�1�����q����Z�eKtd9sv1��*�o�y&agy�m����i.�Et���C�7.w�{^q���&�H��)*0b��ز���#�7��8�oҊ�`A��lB?������"X	�,%qz?������s\��L�`t�f���i�B�$��Ŏ�� ᤈO��t�B'�iK�j��j@n��&�R����hNE /�*��#SP�3N�˒ ��x�nµ$\p���e�GP�W�፿��w�����#l�v���#��첼[Q'vV#
?��D`����������$)��0��,�Cy��١HJ�u�r�Ղ�S�)���۟+���mld���GJe�<�Ir�lN�|�R����؞�k�mr��>`	�9�Ɖ��D�t���i=�[��@oLd���-.F��)�� �'}��A"䏛���U)�ZN���!�h���w���1�*��Υ5��!X�3~�+��Ԉ�H��� �\/f5y��<��|܊���@�7�����8�՞�ҝiB����A�0�/%
V����ŪJk��5�疫�N+V��J��讔��|_<��fZtֶ||S,ϟ��m�6�nzYn�h	@�:��&�D+��@���	0�1�N17jp����#�,W)��{���:���9��Er=@�>
s?M4�'��W������LP���<��i1�f�]>3�� ۔�e\)Vq!c�[_��@�b��N���f�5���� a�����O|��g���e��y�۾6��"���Vp�"���W�˚ ���N�\UW���9�ju�tf*��:> ���Wv�5B�:�N��IϠ��D��o��W�i?����J���{#�e���k/*W3���Bq���$��=�*�1�G'�j�[ ����@g���|�U��'Hc8��cu�
�&"� ¢$mՉ�,1��d�Kf����ݒ�c��p�\�b2fI�3����A��5��8GFG���;���9���Z@�@ļ�r�+��si�0��{8ǛK� #e�����r�{�M*�������m)��G����ZH�)�wi��0��RP7�ʖ�������<�C�X��Ov@Ȩ�2~�fҥ�]�v�	��(G��Z���G�m���S���?��Y9�MQ�e�Y�b*�Q��L�p�J���=ہ������ڶ��gx�_��iM3,÷ڋr�9n��)�f�����lk���`�n3��8���6,hTv�r1/��(éT�^�M���ט�#�V�S�,-w�!���<>���l���.�N�S�J�zg�[k���B�FZe]y��3������ ���Gѓ��qؑ�n�4|d�ւ���^�cz6iy:�ōjm�pv�2�,8J�B