��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	q�v�Z��\R�w�0xtʎ5x5�������v�7\M�k���%n;c-<�<;�`.���B1�7���[�D�\�A��fIj�)����懋�f�7`_�%�E�i�j��yF���^�s�[wg`}vёp�M�=&d.�ȩ$7l	�$����>&R=�M� N=;5k�B���t��7�@>j�c�� �����<�T�3���:����� ��	'
o 	�����v�E0=�(=S� �:$su��
�T��퐣�nXq�u0�pG%�κ6�t$k�%�,�er���p�����w��6���@����jV8U����3~ݦ�G�nM��D������g���擉}�0��j�j������\9\6
���00��?��#�&�3=�ݾB��T!e�?�I�zEl �+@�_��(��6���H_��C$IO}�j#� pꂪͿV�ԲN��z,�An���kz�|X�zB-,���鋿�A0=S����e��c��	���E�]��Qz�'C���3E]Y�ؗ���#HH�l#ZG�y\��
��`��Fk���q�ۖ�ZB��E�<�c� �w��h㦢i��p	��T� K�mۖ=Y���}*���mp5{���]�*29U@ǅ�l�f���^��G9I��s�fb�ׇόxV�U+Z�v.�T�������'6+3����.���!Sd�8���ߢw|h������ �;���&m���mA�2|�'U�,]������CDo	���y���GnӨW �!�`8�(A�wST�j�C���q�~s�6f�.�#I}pD�Ph��?Jy�0���ME�ALMz�^OQ+��y^�p��j7�	-��:�7��Q�@T΅�x8�,��7׿�%��L�'��=H��g[���ou�Jǋ�f���Q�ʏ�	84�ojM�b g�/��X(4?;E(�ɮA��8|�_tB��k2�=�P��;�PrӼ��;·#�Cl�S��`8��5��p��{���{�%N����9�M�7%�ȞbO�9�`��r\ed�_�n>�*j�)Rr���w6�g��E����V�]�eؗ�:�,B��\bۨ����D�du�:qIN+�`�"[O'cY���Kw�����H=��=:'nsz���>���O�Pk�M��3�������;�7�9�_�$H��U��5iS�^GCG�c_�f:�Ɋ����Y' �S�>���z��v�MzRG�7��Ațz�*/	� fh���Ҳ��/ϐbMg���co&]+Ѵ*Sl�M��kG �f��xs��j�� G��\cϧ��&<`�{��d���k�x�˾���ts�����*��br��l͝f,Cu+_�V�����7�[���2N~�rS�c#yIEN,��˺���d�[�Y��v|ﺯ��˩�H�E����w�׃R�f��=�������.�|�ޛ:|�������}bne��*шw>ʽGz�b����"qp}�\��dK16����=��i��7���/<��ŲIu��@��������O�]>kaD������u�(�탵����� ?$�=�$�������%]@|2�v���l-6cF�)a�ɠ�0��eԃ�G���ˊ>'�{��cm~�&vN�谥\B���a��x���) ��𷕅� �@.���P#՞�r�Ч�cm�ɛd�ҹ������F�y���{�6Fg.��X��"˿nq�5�ӭ���V@���a��NK�v�3; ��.<��Tk�|�Uy={Of=azP9�`Ό%��n�q�׹�I)�O�(R�w���d�Ɍl��@Q��zY��@�����Jph�-��N�����-�I[��LE[7l�(�ƾ�.�Ǡ��)����*Qz�1�>��-L�����Bb�6yY�B;�(H�-����81쯡���4���	�;���2)$r��ُ}] oz�4����ec�����<g�C���/�x�����X ���{�e�8�k�o�u�A����(CQXeY�!+��6��k�wXR� ��/T=�R�����_^�<���3�Z�U�|k�����oϢOJ�T�7��g�k<BD@��Ԝ)t�~�����"��Ø��he�#+��1	�}��[8j��ٔ=-#3`b��[�Ew�A륕Lp������P���@$C�k�V���ʟ7J��\7
h��cX9�-d�!�ޫ��;�1:z'�q�\/�Ɵ;{YP�n*�Hb�
;���r�40��Q���T���.�ߍ=&~�5���ʀ��3���|�|1=�o�8�?�1���&�_ZYcdS�W'�F�D��/��p�W���*�"�<�'���!̲)��H��c��\C�kqly�V� !�$��k0�4�ꟍ��_�1��n�D��w$Tzmm���Zb5�� j�ct�ytrL�l���3�D���QLEz��3�DJ��r�j�d���ݺZp�\T�\1op�2`1�LZ�sg�3�7q��'"r&��D�|Y�z�,����a�ʡ����R�\̋$f�C	�@��&o|��,�.���-s��>j�j�`��N��
�2�7<I�n�H�2��פ����~RΩB�oy���G<Z�Ne�72�d�3�#�$�1=,��{6��EP @�$)*�a��s>��r'.�6]�����ؖ��VW���v\�*]��!U�y6����m;�%����j;�Y���M�\ƫ�؇�VJx�s|eZ���V�[U��ܞ����s���2��N���47"b��~�A��!��ՠ���ҟ��c�y��*_�a��z��N�VJ�3��'��Q����~^���`��/��0:t�%��L����x��pe�x� �Y����5~�܄�ę�D!{
�P���ˁ͝�\��u��5�Kga�(L�v�8sj2�s����>W'�V(���{�'�U��N�r�M��1W��+���ڳk���	1f6��4*�ȧ�q�v�H>Aqk����K�S�i�an�t��j��_d�a�x��܌Qq}�W��7���Y\�X��h�di"W�U�i�썑���xf[0��(V���0F�l�_�~��E�e�Ƙ�UAD��;�WtGK�oEB��*~��Mȏ�4�YO��J�r�.�P�K�>EW�s67ߩC�drq�^_�"Y�*�%��Z�?���3���4�x�������s�M杜���tM�XL�"B�WJ�ϴt�M�6?��B�挳K�J��k�����3�5�r�)»�#�����*�U��AP$~.w��YK�"b����ј�����|�m���t��ymyoI�-���)�Z�����G<�;��\V���4����X���2+�K���A�5r{%��9���++~��yX�$���ͥ(�*�,@��ت�)������
>�q��-����i=v��"�h�v.�E�XȖ��ĕ|CqmS ���;�[�e'��Z]t�)�ϗD��4{au�r�%[��\�!�`��oZ�b��Ʈ4HiO���L�(���忚 'M�:7��l&�u/����G��`��`�w$��٭��G�J �ՠ�$���Ȫs��ق�f�m?�[�I�k��!=&��X���cv�%hH@�.�j1����\#�@3�W�)*�/�ɰ�|�|I{��(���TI%��Z��2�����)�8�1b��<3�*CM�����XR>��� bv�UG����04[���%�M�!cU�]vb�A�A�����Q\�p�t����%�M��T!-�IM�_?=���y�>y�]�|Ovg�LhZ+2䦙�'�B*V�VK�����͓��3�k'$A�"|��p�����A؝�%�����4M`¿�w����ɘ�vX�i�� �:W5ӿ���wX{�+_���T��$i����v��hM���.i�?�������4m��8�z�A^
��ٷ�63yҶ{��vk:�~/����/��~S�k4w3�T��P�Q ��]2)�y'%��V=��L�����R��t6��1˘��S��_О�k�_�1V� )��fm{�ei䔚�>i�liu���܍�EX������!�G~,�*�r��>P9[�YEJq�����6$ppރ�4��t�.X\zEٞ�X�F�����iA]C��P�x�J��"����^[�g&9(�ێ���L�y�����<H���c����vX�ѭ^R'���R��X�%���-x�����O,��3���?�&j8g"�k�P�!8qb#~`:�@�I�d�5G�KXR*
- ���rB�ߔV�2G�&��KQ�|	}�8)lz�fS���љV��YF�3x?m�n��[�]Ƭ�=C�I%��]J÷��)ad��I��0o��2���|E��7?�W<�<��g+gx!�y�,:OϽ�*�r���i}:��翚�7(����觿�����b<��`�o��{��s�B�9/�����7���rB}鈾)+�/ξ:��-��O
e}�uq�� !e�����4��TN[�QX���OE0�P�%y YdI��X��j�!��=!��[��/ɚ殘ݘz�+�۔4��}���1]�`v�|���:ƣ��be����Q������&�A��;��:_9e϶�H����g)�V7�8��v��S���������h5.��f��G���`�*�S�z���@�d��� ���
�OIu���t4VcQ����V�4��wW�[YIMk����?dA}�s�m���Y��_s���2�H��_$u���1��Zs;q� ��8��/�L�ϣ�'H�T�FG�5�w��YQ�,6��(b�O�a/��nI�B��'	L�U���:�)s�BӠ]v��<yG����pe�v-�ۻ�f�wn���b��T�z�I�P�j�˸���ߺ|���S{A�/"�0�3]��~�.��BJ1P� �%`��'4�[�I�x��'�Ƈ������:�� q)'���i�9����w80{h*I�f �1~����-�+ {Ә��vF�����P��4�Ky^_�=_u�h�TS��ő��(ǻ%lɧ������	N���XJ�zWŔ�7�l-ž�x�zN�;C��a��M2�pEst�Z�|�|}��^[�r��߼m!���,���T��b��wS��1|0��p���R~���,m�k����Zy�7�$!�M�H�q#�Z�-��M�Ru���>��:H�F����*6���t?AUy��ҷ�(�^��QY�sk��:�	W���� Zr�,vyC�vC���hɣ�p�i���Q�3����jh�;[0��*�rU���!*/�X*3�+m�e�7�[��h�q&i�s���3]�2�p���B �u��Ji����tz�%��d��J���g��d�V(�5Y�g&�!p���=��4�B��v����Ǌ؏fź�z��#83÷a�9���9H+h��;ͷ���o�B�fUV���ց������^-��EZɰ'�&okh:�fk�n�4��0��7ɽs=ذ��bd�\��xߏS�"b�;�G29��é7N"��	�}���S��~�r�c�������]�F,0�.A|�J���4Fa�����$�*%�ꏁ�ch�c���	g�Q�%���ܻ���_%Fs�����@M��C6���*Aޡ҅��Iq�M����1fI:�KhPtnzC睹���.P.~a�WP�
�м{�o��"���F�rCSŶ�������:�$�[�$4�'�C�9�Z�7�g^�a>C��i3�{�3:����~�vG���G��ď���4ƺ�y2�:8*�N/|Ĭ !WL�x���\���v����Ir�g��l �,�"2V5l��2�\��W��[8[~	���-kA�4c?����vv[&�=�fi�}A�9���m�/+�^Z�[�q�-��_�F^�$"��,s�_�%���[F)��"F	��h�E��ީZ4�������)��}�>�L�������8v�;Bj�H?�6j��m�Gd��^^܏��y��!4����������5$��NgZ�n�f1yŚG6�y9�=}OSD�����'0u�p;���f���:��7�nԸ�'��-��Y�HN^m��e]��f��̌��(��`~�K���7��߭,��ށ��]�"����XǏ`��j�g��?�;G�=x����N�>�3��s;��DӯqqJ��,[�v���*�a���:--ș'���3#�	 E�3? nM �G���t��#��<��2�T��ם�ıX��L���V^,��)�����o��g��a/��V�%+J��\���(��(i�Aj
f��/5iE��]&�a3��@`��=������u%���FC�I���� ���Թ�&��V	�m�.�v	�s#G{m�k�Ǣܛ0\Y�]��
_�
?��Ho^m|��6�����殱$]��� ��A�\ke��i�z�5q�6�^HB 4��図kr(�p:�Mijz@X��V���IK���0�x�������׷�d'r\Y��EE�0E~An�u���Ֆ��|�}��JO(��r��N7�T����ެ?��Z.͸dT�D��aN�a������^#I�������5G��\�pSC<�w�H�e.2�(�"��[O�}�JdN�ڗ�1n���^c�#�'�n,�]ؚ����{CᏀq1p��I�L,DHgZ'~r�E�Pq:H�sՃ�Ud$�˞��,�`���Iw ;�����6	nO���!d��0���:CrΓ�Ab������3��n;���@�A�)}
�����������s�K��ļV](�3����[{Ѕ����ñ�YN͚G�P2�9��r����?�����|)�>!�m�"�, 7�Z׌�6T�f�t�.Z�S�h�b�<T�Y��9���d��8S(y���9�� Q��h9���oC���]膱O�K%��������.��Η \A��� 6��A4���4���
&0���/L�uM%���i��z�X��ǧ��6��ΕZ�i] q�3�w�R�;�k]CS�u��"�LeCh4y��tӶ �ڧ��?5%C�ܢ�D=���іIp��!Ǽ�䮊��@��,�H��8�,��rB��d��g\���4<����� �r��<6�E�6�KbO�G ��͞dS`jX� �~^�вR����a4!59��:���H!ioc}*��U}�I����ϼ�_����8K��U;A� ���6��fYa�\YB$^��Dab'y0��	�+�e�ہM#�b�D�E}�,�)_�#����O��AƠ���32Pt�>=-���	pޮ����ׅ̂y�?5H���')Y$*sEq���,0p��S�����i�v~^�T%UU��<#~4�w��ӑq|�C �ߵEw��u���5�@�!o�F_F�x��e�]H���B��CA ����n��6W,Q��5"�A�'dL�A����'
�o��~�&������	�am�-x�b�I
.}�������?�Wט�*~~,ۦ�NC&e�`0}��ԒC���c�^ˎ��֞�"6ZT�SD[�R��-�U���pC!���H��'���1P���nv
�E�>��U] 6!������k�� ��[�H* "ح+@�q�W/$;c�[h������0N��w��G�SI�g��mk�2�6m{�bH� qQ��k��If'��m��/:�J��၃@����%B5�*g|�@�~��Z t�LF
i1_�XbfB(��35:�wT(D�J�4�]%g��Gx����X���ͪ��C�o*��5�p��:.؅��/�Qz�(��w�T#�J�z���H��z�ro�S ����jo��&�azk[y�%j��|,v�j�:Ǌ�/�oTf&�tS٭�:��aЉ��	�<�l�0�G�RyP�K���,"�$Mg��{"��sa� 9 ��
2�������G/�~��$V�M���������l̃�i�����#�<M�|�W�K�H3BIT�5J��|N ��|%����.'�������ق��=˩��׳���Є'4(d�L���Q��χ�j��B��:�/����L��6pv*�"E��p'P=y�u-[�u�JL��@s�8>+�A5t�=��7a��uq|���Ne7���Jq���r��	S����)���_���SK9*��_�T�"4�����eKڠH2��rj�:�n�'�N�m;*�����+��M^��e��&�&{\u����f�J	�n��>�yq~��b�ӰP�i��Y&m����!vG:�z���qBǾ�q�<��ƣ�֞�\"1�A?�-z�*�}�J� ߘ�������=@�(���� ����Ϡ ��Z6���g1�>cT10����D�J=��q�J��E���pX��]��e�����G�'����ܾ��<���:s����"�gl�p� �#��l�jӘ�Q[���`��� v�Js]�&Y��s#6(
9�
�ϝ@�1)������3J];T��#�qK�'iD%Q��k_����(��Z�q�ڞ҇n���c�ͮ ��A)��U�y�Q��^��������'�1��-���	Lγ��*�w�=�!>��"20pAg� at�
6aoBO���8�b�u&��#�NA�$=���|�	��Kbq�a[<�	w� (I81����"�,t>ĳS��x�Ց7x�]���%W�wd�ZJ��fM����Hp�Y�5u��4-���~�:�PX�eW���00S�O*%��29IC���$mo�{�Vwf2.���)�)R�+���1���Ø܈G��^�1��U�R�$��A=�0�q�%dLٖ5.~�UNT��5ǆ��F2��8��S�@��E���O��2m�?��U-8�"�����v$W��V*�U/rE�x�VN�1�>��E �_�~,h��6������ h�%���.�����@�Xj7��뮌)�P\�K
AY@���n�G^�[E9R�]f>���0��F�ۘTu�-RJ��;y�S��ǱD>!��S�+'�@/j �W����D�#A��I0�3�� t��_�α����G��������0ؑ��A] �}z����#��д3�]O�!_���1�
�f�#���
aR�`rJ��]/l��=7 �tlR,&���S�˘�$������JF����q4��A(��w���bǃ��U� ���QM�Ĝ�r����D��s��K�5[ A���Qd���[�]h�ʿP�,ߛ�&ۼbqv+c=L�[�Խ�_�U)Ŵ�5n�'޴���ϗ�y��8�Ȥډ���;{Ni�:q������2�6%*�z�'�-��uGU41���瞂3v 	���C�̗b&�A3Ŷ(�!\�چE��{�-����x�.�K�D�>��03�F}+xr�黝��3��jL��4���;����vd�R�*�O���(�� �Ij�Gp�s���vs�k5�71�k��?|�^��0����GR�\��wi�NSހ�[uB3Ň>�������[�Ad�1��l��~�ż�TcЍ�i>[q��_¤�1'/2��Bjv�֖���l��rgB���~˨-zm U!�P����.�7lS�0�3I���͆��GV����*�
��D���%�|�b&���=zY
%[$���4%AT��/�(V���.S��i^r�`��v�����b!֌(n|��U�yڙ4�.X�C V���{$9D�+Dk+����i��<~�r]�5��k�s�	������� ��S���L$�a/M,5bZ&+˴b��<����3!��̣��&��,J"=�"��ְY��ʈz�����y�F�����]ֈ��̔����{���wJ����ҳ��<;��[3��� ��� ˳s<:���_e��&�PV�J*�_�)Vt�ZMR���y�������ϳ��r�q�����x꼩BՏ�6JU�-f .u�2�T�������w��8�c<��7<"����}�=U-F��e���o�"�ˌȥ�,{��r�h0 |�5r(h~��-�u��W I�a����O�����S����P��Q�rp9�4`��eǥ>{�X�VK����v����9;Qd��qtôx�P؆�����1\h4`ki;d���}��H�BhY�8�J��1�	3�ۣro��$��5�o��Z_��A1�c 9b����C"�1��n�Ұ^�&�+�p)�^�w��vfєM<j��n{tq��lC�i]=��ƽ�P�&��a;�A;/��rx6JI�
1�Ƥ���a�j�7��҈�T!��}�=↢ k����x}�'	VEf���]Η$�¶�t���*����w�K�\;�g���ui��M �vWvB���=IY�
ʖ]�f��4LA�Bȧ�E�p82��X���T<I9�t�fц���ir�~Y_EO8#0�a��5����
X"+o:��Sp+�3!o��4�4b�Y���h�wg@?4�z��Ԣ�$-��*���,A���D��7�6�̉�����U�h�LS�_���(�S��ǔ�O�T�P�<�����q��0���݆����Ǽ�y*�A4��#���&�7Om��g+�_y?W��J%��E�E���.X��v��#�gcض-uV���_���sp���
�Ŧ@-���BDF�d�TuE�v~
7f|ȡ-��@Sw�.�4��.~P�GW��%��������ؐ���4�f�brPj`�Ș#L*@Lbw弢l��V����A8�m����#�@P���6��>�Zkq����i-�� 0%�Nr-aӥ�j����;�c���q��R�}�p#>I+;Y5T�\�E�L���9�hJ?��Y���;���"�ĭ���K�0�L��I�t�ŽqPzp�A�*��� ��W�y;��1�h>L9��a)Й-0��VS���'2��kM��u�Z!A~�L�C���X�;Hl>���^�����=��e����N`�&-N�.#���,��@��t@�ٜy���Ѩo���b���hDya�Q�#f��W���w����=��8�5��Ȝ�r�eY��pat��Y���a�ߗ� !`���5<(G�T�|t?�r����FG
��!5\����S�t��(��	���k��g^��!ͨ)PY��@�e�h�n��!���+���5�Y��C�ō�Ӌ[3�Ίe��y�4T���y`d�i�۪R��-�E)m��!��/��Dx���^��W��4$L:���׈Z<�*�Q\_�z̙�9c�1J���Z��V�Ӝud��L<�A�UqZ����E?�)S������Ѣ�ID`(� ��CH������l��4�����q��@�B@�����k��̵r�1ŷ)I�r����z��d��GU��Vg_"�5����R��C�|1o��7_��L3��\�d7�y�S�ŭ�&+�7?�k���; �ۄnFP�^�_;J�g�
D9�mo�DV�Cf��cG��Y��^߄Ut������q@	�]0Z[����~À�r"6EV9AI^�¿ω��MɋZ �3A ��qA�eN��et������Aq��t݁P�:F��ۨ��4�ܗj'���4#��N4vJ.�~'ށ���5C3]]�W*M�|>F|I��y��-<�^VN�qSz%0�v����=��}x��[����
]Ѳ�yI�gYO���)Ȳ@��Չ��I�檮9����7��j��	�7x����o^�XbIA�������oľ�e��uR�{��^�U���c�{=q-���X�Q{F!�KKR`��x�I3� P=*#m�����#����ກ3������^-9�i��>�A�\Z^[��9�g� �Zń��O⣎�1��9��') �}�����jo��������O�6>j���Rǟ?O�ܹ�j�����Ⱦ|oږz�u\q�� ���9��H  ��q��Oe���O!?u?^�"z$0���\4S����Rt� ��w��k]�Ҽɚp��!b������-5��������
��ҿb��:��Rx�*�/<����ɫ!�&ʕ[��ueuU�@SזY/�� ����-����qs�f^ kM�YEuGT\����W,qśGZ�X|����\���J(ǟ��sz������7Ҹ�/=S�n��3(�[.W�F��V��q�N��:��W�N���i0�c�w�rzC+i��ꟽ�]esй�8�$Q�{s�\�K��@���@�2�� 0Pc�G<}X`����7��n�f��:jPn��IO��:g:��+v�*��+EZ˓�R��|�ڵ�V6#/XŇ�M1��Z�����ڻ�o#��Y��~�g�$�<@N��W���)���I>��-���\���}��q$sU����=OS{"�������3�M`f��f&"���\�����/���GF���U� �b���*�H��ut��n�U	�|��B��� ���-�*�'.�Al��0��������-�elL\JA������t�|���/������Z�ɾ��r�sx�`�������1#�Sj��0��~I6FR*{����7������N�Rn9�9�[p�0N��l!�D��	[4�蘉	+��MK��U��ḡ*p�X �3�f� (�0"�l8f.0|����]�����fhͪ�����	@A��X�Nk!�����-�q�vĶt���,�8��qҧ��y��Θ��oֹ�niOIY��ܑ����v;�������+[��`6���"�'b��G?x�r�b�2�$t.��lpy��8D�)SA�S�m(�I��u���c��|ے]����li߃Y���d�m��}�W[Qߏ���jȈ���֙m�II�8�@����I����0c6��3�e�����=�gƅ���=:�~!���<G�GJ
/#�=pe�Q�V: 鮾���nAK���z1~+�_n`�Ws[���#JƖR���ŅlQ�o�82���ލq�`�4���ZY�g5��$M�&�;>�_Es��%�$��f��v�}>�c1Rap.qԃ�H����V�0[�����{7'���@����V�&W�+hd˽85�(�n�1R��3�fC
���	1	km��kB�q18kS��2k<,��K��I� �%�pJ�n���d}�� 4*����A�F�s����޾��m�ihZ��a<�<*����
Xh�$P�BL/���m��Y�S������q�7!M�?}N��8Ƥ�:l������xm3(\(M�5t�:�ҳҎ ̷�Pw���B�`A.�<��x"i�B�'1�E�����*���:jm�G��k$�@�s�[���WZ�'&x���'�8`1R��6���bίg+�%�Z�y-TK��ϲ^���pjʊ6��MG����Ds�B5!�y�n���T+2�aTk�߽���v�b;n*�!�%� ���/4�@�Bo���x�����㬀)&c,<5�XI�OH+y�>��T��*7J��F�΍����@���/|UK�",aU�����Qk���7,c���K.l1�������'�k�F#�eD�����ȝ��5��-65y΢�^���>�(�$!c�¹������zry���N���A΃F"��3���/w�O_Q����DF�u��c�𴾱7z��Y����IN�B�(���	�ˬ������;�&q���a2�Ҝ�襉��6ȉ���rZ�����gŨ.���L(�h�Y����a�o��De�
�qx��9ƍ�
k{6'l~��l��gp�Ȟ�v��MƁ)�MR*�-:���<>�����g?/Y0~.u:�y}O��v8����b�	���E�B�2SVD^��DQiV����x��\��d�Ś�ܷ�xgYb ������q�ogH�/NO!��O�K���_1��D��ߗ���g���CVf욻��A}�
�s���Sk�Pӝ��R4J���S��Va\Q�k��%��g�b��\�=�`[���5N6(�[\�P��8��U$��|��V!��7��MQV�K��A҉������g�%;�V3"v�UT��*&l�³N`����xHU�
�xj��֘��4�C�%��$X����z-]#5.�:A{)�>ĭhH�DEzj���W&c���sR��%lH��}7�asiR�l-`���/{��%�����y盄4%����2d_`��7N�gK�.k�u��"�2�
�:!�4*�'�ɾ��+�8����>x��`�i�%˖'d�s�i2� ��]��`?��+��t
Z�`���8�Y�#��1�n��\-k�?r��ekd���v��A%qU��-h';�q>K�vrJ�b��Z]m�+v�l;4���0L]h�ޓ�7����hT�{��q�&�V�!�$�͛cQ·J��#tM�y̪�5�`ċD��h���e9��|��x��X�X�N���c{@ǥ!����h�.M��f��G��?x�w�$����{�xt��M�Ԍ�I<�T���io[q锋B��JҺ�.s.V�ٖ�[]9ڻ��5�հ�:�;=�`���"kLk�*
��S�݊��u����a0�u"���Q��WT���-2EϩsE�LݹnIc�-��<]R#\	��ܔ�e��b����ʡ���!�� �|�$��[���BgS[�e=� ��r����
����"��TY���Ex��vP�R�j�*���?�KF�IkuG~5��m�!'�^�L7Շ�5�-j��^�5K��0��p#����P�B��:JA�5��c<D�a��A_�X�]ސ,z�T�,����І�vɷG�n�8������X�)�B�T� ��
�4+G]Ț�|��iX���^��)����ǂ�9�ko�a�,��SNeBFi�HR��ߖUCC?��[h���2�9�OtP�`�Qt����hc��d�m��c�IF�&�SæB�F����[�3���`p�I8�=6o6���{�<'M*��1���E�Ge<�,�WjeD�����X�g�p��B�'��Z`�ֵ�HߑO.��Yq���l���gXd��Ǌa�x_b��߼ԱP������T�M��6��cs�HeX��jμ;1��&g�VME��.儮v(aE�#���T�h�ҏ"]����4\��B�F@�f�N������#^��9�h�F�I〮���S�l+��["xl�Ou�՜W����`
��BX]�p:�Ƿ�=4QRIǨ�x���e6֦
G��uJ��h��7�g�i��yYE7�d�zb@�|4�I���b��1�<:Z�VC�C��Ȱ�5>��5D��G������*!����Aۧb�9M��#�w��TX�L��E�r-NJ���h�KN��s�/�xN���B�f$�b� ����6�]��R\*b� �z����Lˬ�Q���N�%B&Tn3��H4�ݽ��)�#�j�f=s���yB|��-�L4eS�i��h� �uEB�����
Ǹ���s���|2��������v@�c�9`7Ïvv��� `0���n\ص$� ���S�JX(�����s�q��_#�����;n_�'S�����&�ݤ����j�^��ڎ" �/y��D���>_���1�/�K�-��q���4ف���1��kEN�>3��8~�\�i��L�Ǒ���J�;�ي�g�9��!��8������F���2��	ZRb6��8�1M�"��c�m�F���fl2��Zm�-��"9�q�V4X��E�2��~d�ia�p>�
H�D�
F��2���o�:ڊؖ���wK�pꁤ3����G�Z��zyH�7��!P!
!<��u�Qz�_��F�E踵iH��9°W.��p�lx�f�(���Ɵ�4Q���V��+���d�p̪[Zsj������4a�&b2=�<*���	���&y���Ɯqp�U4���� ��� I�h}R�����������@7*��h!&�Q�d��T`.���V�,@z/���p�-7��j^Mp�9��y�H�]�@i���I�O���/[SZ��i�}����C+W�E��q�خ�KLܳ�~1�0R(D�N6�g]4����DuG�������n�2��O��b�������$�B[�����	��V#Z/����W��F,*��=0����a��PD%�C<�`}���!�m�Q��D��-�����sŋ�0{�^>Z���iR������1��iX�qul�&�
����Q8��;���}�_�(��C@Pkv|�o��Mh��
�(�T��u��FG�2 )D5�-o�R�y܊���BѨh�U��U��F8�]������H����?�,�����E�C>(ۿ7��Γ����,��nw,�4�����]��־�TNjv�:�B�[�z���[.�gCc�t}�8���}��b��uD� Z������;3P�FE�B��i���I�	�<Ft�?M���葈�4Nk�:g�=���K%;���"�:{���\_�[���]pȅ�����0��=�����8^�e�<Z�@�xB�EO�Iug}�B0�ܾ�{�����8������V���K�J��%��=��FoZ9҄C�c[*q,ű��Gwӭ��`�t潳�?'	��v��n�L��Orp1��W�X��D��Y��c�����jP���d�)DԊ�L�9�0�(����2���Yt��q:	�2�G��Y@�e�V�`v��D����G~��-���"��̦8��>� �ݚD�c4OdiH�7V���^`�H0
� +�7_{�쮪��-����zӢ���)9�a�u8���4����'g�S�}��j�i
5x�D�x�&#8���~��a�X�#��n�N���!�@p��|�#-���ft8�J���1��x6D{}�s��wB=��G�] �2��H� _��Ґ�7��H�7;��j� ���@��_��4�}XNͅ\Y�ѝ��5��e��foRt�5hw42&eϾ�r�8�w�Z[9��é��V�\>+�	�~�e\A,��!��.���'�&Dc�'> -��XE�yسhuW6O�|��Z7zd�۷���bQ�iU1�t�oy�� x+(���-E�L!�տu��:v;�'����B�Xu������{�>�87��
��ިcRER�OV�l�Qm�������פ�n��*��?D�cYaU�Y�.�o�;.����jP�f�V\Us��}��hpx�D��C�:��Q�>θZ޸K�r��D�b7�O����ߵ�MCu��]˰��.K;X��2���g���f#�9��Uj�ǚ:�$���?9��`����Z̜��J�퐠J�>��\������zB�v�h�/�KV_%0��P�I�%[[	欯�U@��HTY ��A����NcuT�U֑����삱��1��.��EHG�NETDK+HSP�/�)�I�?1B�{8�@̈́���09Y��(l����^��/�>��Z����r����Z�S_�&Dj�;���u`MA�w�]��vɞ�1��*��fj�s��[����`����~�]��o"|�75��8_1D�rD,�֗p	�48����r6�6�G+)d�^W�������~�j2�P�Gm�����lX�0�p#�T�&�m��"�ݍ骙ܲ���R�=0u�n<@JLHj���z���aW�!dzڷ��� ��bo��W���q���NV�>�<�%n��+W;�SV(��](gvK4�� M��+�&�I�/��H�Ʉ��s߅����]�W�r%Yx=�,k���b�8�l!��XF����$.ɹ�F䦘Uԣ�&B
bY���f� �KgOEh��a	*'� �|,���V���yY�1�N4�=� �ߗӨxB�8�pé�,2���6�܃h��`�sv�B�N��i$�ؕm����Y�Γ�=N�?o��]�m�1N�Z��˰X!�֢?�Z�c&"Z�TU�u?-����zfӌ���dJm�K����\;�a9h����~bW�#��C)B@�9�7��z���AU�mN���sȑCzo���,*��j6d��d;"����x����ZxC��8��'�pŖDcnq�F��6�s���7�(�~պ�s;�m��`D��`�2�s�/8�+U�Q�n����s���s��D�^>��)l͔$h��x�GAO~w+����(2��k-�$�
��&���&P$#���;�ѧ�����|��⇩�S������b[�f`a�h�f�l��W��Ig��T�U��;A���<��ut�G	�9A��C��_a01�jO��$�YΎ�AQʛe���LC��?]P��w��v��s��e:g���B�7� �7����c}�؝YWԗ���bZ�I?�;���;�������x��\�1<u��y�@#��R��lZ�~jXq��\�c���qDW��՟�i�=��m���ܿ�i�Wb�c���r�����H)ƅ�l�X�&�����-{��z+�F���l&�*RY����E�O.V] �����mTY�(�q�p�5dBe�ce����bź�9ez����x����Ѱl�f������[�:����!��$� �4Z�b�U~��	,R��\A��'h�s@䕯���W�ieּA%��1�q�w���$�#;��fC��7�H���$�qx�-��jq�%}�H����;��>S��1Ao]��A�v*��ˢ�v�f�����~���+���-׎���� �Y}��n��M�C}�#��x5�y	��o�ȹ~|�P�L�r��tXIb�u�]���u]�$����Nfٰ��*�c#Tbt�|W'm��H\]�V2D���������]]��X�@F�eٯ$��Tz@�S�,�Ȁ�D8���mUE��Ihvt��o�]��'���o�(/a�譲����*�_��FɆ^����w�X?�:GS��X[�d\`D�Q���&����D��f����"t���:�s*�$�e4ɰe��c(i
t�[@�F�V�ACS?n,���?���(V!�9���&YT�c�w��lZqV����rT|�� �fw���M�a;.�Je�3͜�{䶩X)~	+{�;�-�a���ڍlG��A��q/���D8hc֭yv "
� ��*�S{�hq|6�:Qx�H�����H!lQ�v�=��L��k�u>SC��rOvk$0�Q�A��Ϋ ֽ�w���;8��m�b/j�8U@��w��%��z:�3t�A���C��+_����)��$�[��nsF�K���A��;v�\?��u��`�,O�5����z@�+������|��@W��qA<ð�˄<h��?�`��n�]�p@��:b?����������u����#0swI@a3����D�=�C�su���l�r�IQ��^��՝����4�P
"�^���V{�o��$��G>÷���ݗ�)����ح�M�#�&��:�������]�*���d��7���:I�9&@(��}��|/P
?�F}W��/�������ڻ����"��p�&x\���ǒ8C�	�mہ��~�a�sZOQi����w�X��)��� "twz�4�ا��� �;D�{"W
���|�]���Q�K���q$돸ފ��_*����yBi���hd�oE�/]U�R�sb���k��z��*�ʴ3�Wa�0�,�;���-�X(�'�j���"�r�m[Cj���W8�P���XU၌��|��ec��ǽ40��/V۝}\�~�N�*�;��Dr���"�^A�}Zp�܃��p�X7仉Ң<��6��H��X0�3�$e���D����,�{GҨ����A��`��H�GT ����c��n�j3�q0-&���Wud<�V��-��I�5��\#'��Mk��
��W�ˢ�s̫ڬ��~`�G�C����~�����XG����σ)�\�q�����S'���/��0۞�y�;I{��'>t<~K���*Qh}	`��*��َ��YO�=!�efU�
T; #r���</L�6u������~I`�-�5H�G9VN�D�(�����x22��P��άզ�s.���D\��W�"����4�ʋx�f���|�������!a�/����L)��0�a����ÄZ@��N�h���Ɯ:���`�G�\!gv�BV�0�H�%b�U�gb��_JHq�U��!�WK�s�������0��Yu�W��㎣�Ƅ<a�5*�m���-�g�Kv�	m|�ɉ����κ
$���3���l2���鐹o�<�h
��W�'�T.�2���VYӋ���GTN� g���1VoV2D�Jc���ѻZ�k@äʴ�sҚ�I�ܐB�B���z��F�/�+�֊�
Wb;�����a���4��{I��̄U������T*� kԌХt�\;fzt2 ����̺gl�E�H;4��NV�Г��
^��;s~~��+�g� ��3y��>���B�?oR��3W|�Pۚ(V��[�p�s�p�kV��Y�Kz�@��w�H�<��l>M�Gw!��t2X�f�SXC��7}v���Q���u�>G��K�G������ؖW�he��ft����R!a���#�I�6
�&�t&pag^7�~X�1�T�^��9ƅ$�K[�ֽ�w<��ߢ�18���	|��%�{���7��Hݴ�9']襄Y��lG�&E���t���{9��l���?z�ǓaO��0i��k=�D^Ĕd3�fE��(�C˾!!��� ���9X4+�ݶ��}Y��E�����\t|����A���ֽ8=��7F���x�<v�pЏ)w���+Q��= ��_�Ս'�D8f�O
���^Th`�wQ��-��׌�̲��Y�P{9W*b���syǈҔ`#;��+Ra �j�����
����=��8X�����eHf�	���]@�TQ�s]�߾ɢV�&n1�oa�+�.����B&^(���9^n���n8�Ub��L��A�M�E��U���
=1 ��b����m˙56_Ƿ�vT���������"���UYR�<5�`DN�4�\W�6���ڿ���ep��1}������jTIֵWY��&n�W�"=�
gh�J�ܨм���J��Xr�:$=\dZ�	�����dkl��B��ȋd.����S��Q��(X����!�rGI��5Iv���B��Uu2nB������6k�Ѿ�T���Vs���v2Z����ۆv�cHɭį�5�����ȃ�p��䔄��y�,&c��fԬʙ� �4䕴��,�T8����)�4Jq�ch��Z-�����y�9�B���u:�{�f*�S0M�A�.�ރ�ɱq3a�^pC��_�n�fx��չ��������]/C��?��~&�W%)�t���)��W�6���q��1����KN�k�PTR��JA��_J����S@4։n5Cfh�o�w���u��\��m=Q�	h�K&[Mg���8�Q]+Re��{ל'��Ad��(6i�ʟ�N��s���z�C}�m�&�����/\�9�ntӴ/X�Q��`��fc�9 �h0�=J��FZ칟�78[{�\ҍ�7-���aS4y2��e���d�ŷi�A?e��F�5�u��0��)����o�A���~o�8'�Z
]�Q�A��T
�u;�3��FP'N
�o�;|�1��Cd� `ڲ�4��)�6�X�(��T��ۈS-�{
��GC��@*��J�7J���7�q�ΰ����=��.���#x��@P��"��Q�p`m��K�OHe2�>\���.��O4�M�v
�<�?�4���P��� �f#�	�$���v��Os,�����bڔ�}��pKki�8��D�0�8Q'�_\%��Ē�Tj8�����4��J�m�%?��-Z�6��3?��X��u\��.��1�A��j������>:��.�4���p�7���;��s�m��>�i��txB�;���gʣ�+B�2��Cvf��]����X�E�������oye}����B�1Ei�C.��`J#���4<��^% ���V�$����t_.y�'i�ѣ�N?�S�0�S�v)f-�"�D16*��S��:�)*xe����{���1�OwO�<�������/	S��x�؅m�� !Y
��5��}�$,J��D��1�|�^��;Ǝ), �������3��%)i��k�9��ڌ�޵6��,l��A�w�_T"UwS��z_�Ζ:�w|�b9F���{�.F
B�'Mr�����$ ��[�Ǎ�w��w zC�k��{GV�V����vp��B�������܊��a5�:�w�$�6#Q��� ����)�w�?B��~��&Jn����n��x�&շ�}��\��1��drќ������5��wh���p��&pd!��U�;���ؕHкO���->U�d.d�����U&��}d�ߴ3�g��-}�W>~�	���~Z��B`��	k��+���s�֍Q�g۬�_��#��H��c��|�A��&�߰%h�4�S��>Q.���|`~;���RQD�aϵ�<�x�ݕSH�q�！�]�F��[��
�����J��B�,�Ś�h���˛7�֒Dᓌ�P�̪
Fr���'<=x���U���3'���K��飑V����
<���@*�F8�v*�s��hػS� �r�ĩ�D��nڬ�a� �1�D�2^B7A�Y��"��Ɛ��`�0��5}ߎ�0^������U+�?�0hǉ�P�Ve�,�1б�Y���qwKN��V&�*�4tQ�E��\Bϥ�����A����[�2�����0��l���H{ރnA�]���G��:h���NB�M{��,�w�cRV��,@��(!�&qA�?��aG��b�_�,���i�)�@��z�=�J8���UX�u�����/�M�>�]����SYX�������\�@^	���ľuN����Z&�4��̻�K��K�������%��i�;[��P�[��{<�(�P��������G�=���yh�����)�y:�j�4a��G����8�U���k�=i�/v�
�6�jBG61�T�}7|5myqή�@�_��󞔁�����EP�)���jH�U+�0�c�s�ů@�� <U%�Lԉ{Z��q�m�f�7{�B� �FY���ޢj~%�/�T>�^p��t����%���u��*��kސ�6�^��taX��m"�_�?��]�05i��QK�!^�*����JqlX��6����vp�Yk4�
~��O�T���u��Z\��D���oo���ڨ</�/�>�����&S$��(��й�<�AU�@�㛙�?��iE��оͰFXH��R8��a����k���_��_�'ss��&xФ�V�ٰt��?��|i�a^���}���	��νׄv�-'��`Uv����V�z���P��3CTp����k�**��e|k�?��ݖ`:���I0�]����ݬ�}��ꧨ�MB���8H�-�XTP�Ԙc�z���m�l7�5�iR�|���|K�~$b"~HҡiMw)FL.�N�+�r���-mܑd�ǜ�礮a� �ש,R����I�=��������HW�_��<ލ�x�w��p|m�H1��Yz3�ٱM�{� �_>�qj��o��Jid����R���u��=�c?�V�^����Mnk�p����J]UH�j6�χ�%3�41�7s�P�2��UzF��lf��/q�ܗie �0�5y��k�rP��)��Nqxt褂���^�5�.c�l�b�����oG�����;���͢8�Ȓ,z�6��n~�o��B4
R;�2x��%�� ������0�����]��v��r�E
:�3����I��-�zMwX?��汕�Ɣ(r��Ƃ�Ь[G@�Br�<�K�/��4���<k�o�-���A)�C7 rm�����~,@3!f�3yZ�,���"P�������O���_��:##0 vS���6{HD�bo
Vk#��}F�PR��*����y�4��i�Vl���/\�J�0�vP&t�n9»}e/�~9�����l�wm<��#0�.2���OJ�ŮPzaN��lɆ�w������&Y\4>����6���+?ej�RC1޾̵����"�E��b������`o�.ǟ��a�U�sq ��%S�b	�h��S�a��s�d���R2�+6,!�F��0��ۤ5�<�?��e��`�P��7�]"��%b����V�������K�H�u�v�~�H�@��@)r���9�N�Q_�W�W���W��]���1T��)��UT}��X(b�?��V{O�]����P�w�~���	�ϟXѠYL�t6A-_�|?\Y�A��' �d`L\�:ο���:�UQu�08���o(XI�zV�A���MO2��!�rxo�@�UP�d}c�%nM�e�C��<h�4R�8�4��P�3�Z��:$(�<�H��Lq�L`1K�ȟ��<�'$�YZ}@�s��l��8Ō��&�Q��jS�t�g�,s7S}
�U�H:�ѕ��5t2�߈{���66c�"D�����F\,�).�v��B��':S+��@a��r���w��1@5��]n�Ș~^���|� �oxH7���\���5� uw����	�x��?��C!�/���`��b5��IlLT�*�0�$��Y�\���7��?�/p�!�q�`{f��EE�:�J�E?�(n��W<�h)	�#!�jTC��#p���+l����݊�v�sڈ��+D?�sx��c�ZO%�6�+箲�v�w���/�d���[o�1��V2��&�D�k�ơ��#�Ea�;��c�U��-������ ���Î�����ys�c�J���j]I���q'�Sģ���S��Z� /E�uX$����+;�TQ�[�i��;�8�_Z�t��9�>р~�	�-��[ދΨ�kIk�y��H�bҸ<@����4ve�H��+����I,Dq�T ��' K��� -�.����$ʭup�=�E$z1��_�J;����Qe�V4���8�S"����	Ǒ_��UT90s.��*h$�O�~bXR4=��!R���j*)��oF�#���y w~�0�k��.Z�bl�Í�t���@���~��FէVR���;���so�F�����������2Z�=�9OX�W��Bť-a~V���0���J�9�&���'8%�&��{}3�q@��z�������L|��O��r��Z�f���?���[��6g�ܔ�)�X�d>Z��$ ��;���������!��k��}�w�̒��K�?�+H�aB�y�A�iU�"��FG"��nCl,.j�+왣���=�Z�1|X�7����j99 e�G{���ߛVnj��-j|�Z��'� ���|����%ݼb<����g\�,�/k��߃����_ZhP�ܗX�j�����}�Kڡ�Puy��~)��Ta8.@�i��ۺ�;5fA�2�Mx��k5��M�Y��}�G�B�or���x/[�Fݏ}�,�;�(a��\ҙ�[t�͸)�}
�l\e(n�v׮�^,|�z���;�/.�$�X2�δ�%�'��m��fҵܦ�;��f8'i������<)�&�l��%Z�T��'��Ң��~�;�Um�Xo�<'�9Oj���/�au����r�
�#�
.�~�g�#x�U���C*
Y�軑����F%�.X����'&}t��,S}��eP�'��r�y�Y����lbo͖���������L���%Ćw�Z�JoBÓk�0�R�2�h�^* �7އ"f���<m����`���D\���Xҝ�(oi��|ޔ 3�UԄsD���5BKnñJ�si�R���o�aٞ�K��%��������zo՚��*����1�u����,��=,�b#E6��j���AN&�E�P1��i�A��W�6~�;n�p��c(�V�!X�֦Y�W<f�8�@K �/��X�/��$��r*�J�ʇ����9Q�f0haebNZ>_�D��0��'�Jb\�8�M,��}�Dߤ�Ȓ�e���nܝښ//*�����~tI��碄�Pj*Va�N�Q6|��8��Nd8#�Tc�<��� �p`^+���s\�F����>�����98m�8t���@B7�f�ւM�њ= ^���-s��]Rʻ�-<�UqU�d�Pc��P!��]s���g��4`�\��fW|��R�vb��q!�؎�s�{��0�i6�K���I�J��`�k�����59bs8��Р�4Dc�ki��]*���"Gǆ�l%΀~K�d���[�������i�� ����xo�3������;'S�='��j����"��hBQ����;����S��2<�\n{�G�2�!u�K�������&��b�p�.
��o��B��b����F�)Yuea4�д���(:]u;>\iA��=|n���#&����I�Y�7�S�|/�	�ݖΫz����jd_	��R�qW�j?{,��~���5M�(����rV:��٥���""��n-"n��.?�?#�����nF���l4�\�@����%�NU{�!⺛��#[��W0u(e�J��=B�E��:L���h��G��O��@�+]�AQ�Á����NYj�T��n3n? R�`	�����T1��2LJ�cq�Y�<����M�ǘ�w$y'.�c��t�~��/>;�)��+k���/.B���P�,�+�3�@{PqW(��g)�|�+ݬ�}�R 1JH�5ʥ�W@��۷b�5�����@�7��	�O\F��UPiS�[�לH�*'�ߟ�t��?����\�=�XqM]y�>V�w?����-�(	����d-Uu$�W�#ݓ�zI�`�ٕκg���g(j�J�f���S��=��TP��{���`+��Z㒍J�<D����[��_�2�X�ȧ(ۮ�:�lNG��MƝXX��-{�L�2<��x5�a� L�����֔.ͺh,�%e�����
�gp&��R�ٖ(W�W�B�1�d+�]|��b��S�2+�'�"��Ng��Ko�����s�����`�1��Lvr�ښ��b=��&��i��h1I]s�փ����W���5 ����i*7-�M;ݕ=�3Z��0�>ҷ2��eq���
��k<�B�k�m �u#A8��8�kkد�j�H%�íɮM-d"�X�iv��.���F8U�I�:��j�-U��Y��MCp�yM�<�V F����llUb���kĜ�Y��w �3�4�0p�>�jp�X�6��OQ���0pf.��_"������"��T�ʭ>	Qd�G����o$,��*r��:��������Fi�2ﰸqYT����=E8�����L5�M�F~��9:�$�2"���KN����>����ّ��^$@~8=6�=[a���ª`?�2�Q�W�AA7l�E��\�<��ҧ���A%�H��$8�*X��"�4F�J�/�i��6�� ~�sk�QYk15<o!�����m��s��(]e��C���`ݐ��w�˔�,��(�]�'Q@ے���fo3{9�.� >�kA���m�x?��������d���zS?u���y�^�ͭ^�0�uf*�-J��fp'��.��j�
g>�7�?�d�h2���?}T4����Ke�}��8��N���F"��p/����@���/�M�Z�ݣ�|Ξd������0Y�:j�cZc�6M?�l.Ymw$d.Z��SU�0\wk���I4��������y}�=e	I���H!����$
��,�n�;�֢�?g�J��h"�
��)B�		�����mi���V��y�a�d���N3�i�o�i�xl��4�tS�*��ְ�F��m�ɷ�j/�R�L�1i���(���1J_���啁D�B�5c�͌_ea��;���է������k����+L���*n�j�bX�wu�Z.9q?��[�;ܺ�;��D��,g^�%]�U�.��`yy��~�x����ir��v�Ō�=�]uS��[�l�����v����I��� ���pE�N��1b.M��l�`c⽫	l��j#����g���h��8�Xk��`��^�H��)�=_��}�����:y"�B
[pY�<<�9k8�:�^�D(�a_O�9*L�J��<v6E�%b^��ک��	�}�\Vc6`/���BN�.��><m�I(]C��Å�ZJ����� g�n5�s�|�L���F�@��	�|zT*H28D��L�z��;��$)���J��e+ZJtV���u�8�-u[��7P�c>��uD�\�S��*t��c���(A�a}lu3��	��� X�D�`(x�*!%��"ZY����E֌fU���>]�AƤ.��1���O��^/*��t&5eBf��ez��JgM�n��ѕ�۰�	;$iB��(_��c=
2Ҿp������Lf�r�x=G���IWB(�Ǜb.�PD��T�ᰓa�+*�cw$���ӯ-Q�~L��㝧r���Q��[Z��R���.Dƚf)uCR�>�gnO$���B�ݐ ]�5,��@8��Z}E��P
�;�o^�9�!��C�9hq�UF�W��"�u�%�
Gq�����V�*�,@�
�'�"�69cy3���쯊!�1���� t��V?���pѤ�;�$V����bA2:8&���Dɓ ~=��x�c�$�|te�R�ߝ~��l� �7̹Cg'.���b�c�(f&�L���.:����28��OlQ�˵��Qn�ܒ���4��!�\��'��������O�NّR�(�M�KE�����<�k�$s'i�� ��E�p�ܱV!_�e��Y0�1Z�~���C��鷎dc�������\��M�����c=�\�)�C���$�?x34 �r_6 �c�x�ܔ���@M2��-�3'���H�e�z��.z5�d��v��z9�*��y�C��;W����6+���AE���(xj����t��1Db�vu��H+jSgq�0�Jф"E4�!�l��Op%�j�%`��d����O琒[��8�Y�	�J�d�
9����	92(C����|ORw���g��R�lUs��fmp(����v^�P���f@������=*��yp�I�Wy�e����d	o奱�du~�nf��u���uRx�/����xGrT�ЄZ
�^�)���6���K�S*�]/:A86/�d�{K@�0.�f�k8�?�����n��zs�q*�go)�NO\7���Q���v��MX�q�ɚ4��p���
�sҠֆ�Ͽ��^��ˆ��>"��L�j�`~%���ʚ\t�+]��v����)�(��uN�1�.�a�M���Vڲ1����@��oT���
{�ȿi,���W�y��#w�i@��"X�hkJk���vҒ���,JO�5�nE��@%��f���/��S�b��;'�ێ���A��)g��c p&�"�����hN���u�(9f~dAu(�~�#��yDM����O-����}��kg�N�|+]�E�Z��H�{ʐ[�o*�p���a��j��������Q�Y�m�O�D$�'��n�����M ���ֈ��=K"M�%H�i��%۹)�`댏C:����^�7��2�S!W���9�y�o�����
���?S#	�ǤH-�G������^����f�2c�vy�z��\S��C��]C�V{SXt+Ur��fN�$�Ç\�X$�"CW�@���R���5ge14�����(���ۿ�M���A�U��I]��:7��Ah���Y���*�O7��S�G�o���N���G�	��8f�+�[	�`Z�/���N��}ot�j4[m�Q8�!��i=
l��o��9F+"Dn����� ���i:��Mm;�-aH�w�m�JLG|���a��� ��J�GU��f�܂[���_�ظ���b�}%�+�n�5�	_��A˃:���Mg�BsEL�Yp��${b��uB�M$���dAeQ���olGg�?���yA�ȅÒ�n̓]�?��A������.USk�G�u��^m���|���~�,Z\J��?$���NU4p	͓�s���p���e �T`M���Ǉ����)KF�Q�W�?誢��g���}�^(A������B��E��d�K9MizGBX��Dz^cC5�Zϱh�����ũ(�JKw6Z�#���D�c��,�<�n�f�~�BY"(�L	Obe-,����a�*���C_
��H�跐�"tI�1l]2��\l�ϡѢ��&�/�	$L2������u�F��<�NZ����/��U뛽Q�I�b��&��"��'Fo�X,3Q������*���XC?֋�e>h��=��w�Kڎ��o� γ�ɷ��{a|[^>E0 t�2c,+�����O�%�mD��l��d���g������0��u���6���#��k����-���I�ᜫt|�M������öU��o��:��( 9h�W&��F�#���;`�M�,��������L{T5��D��]c/U=q�б8_�(�+?s�D�����=_�P�;����ǹ����b<F�!;A��k<U,D��T�;�����]q�`�HW��~����ii���gs�]�����g �gU�8���	��hcM����22ƄƎ�)BM�J�'t����Az��Jm>{+�^���m�ꗓd$�:͊`^ֈ�	raE�fB�QN%� f;�A�j�9dwq�M_��VT+�pKvY܌�2|<�?%���R�R?�@�ɒ���n��FX;=�q��×~���Mv��Y�"$�/�Kr�=����~��}���~��/Sd��5�3\mI�)\ڰ�%�!R !L�AM��mD�Z��Rb>=)����ǹ��c�N뛪���2Ż�E+0�	+Ùx2ņ���'�趵�UEL��a"���F'C�D��^Z�Ь�8�vLԆ���J��pK�BW�4�SJf�����z�F�P���d� ��P˟G�u�Eڤ�� �}m���[j����5�;e��UE6�埂��\�7�f�����Y_�,Dz3�[�n���̗N�Bp%4c���j����7
edL�E�nh���Z����h�� 8ߣ�0�^���_� ��l�=3�*� �{cB[5\*�L5���J�L�٨��������� =i\ԧ�[�"�J�3*$++MբO���9�R�=�!�	i�+�J؞|�|����l�D�Ԑ�&��, �(�LC򺌴�������{������)L"��QQI�}Il�<	��nR!�cV%~�Nb`N�6hi� �e�v��x%���7�L���pc?-�����	��A�{:��Q��o�o����Tf'��LD&w�d�s�T���)�h�,�9�1��g�����-W͋lH����s��c�FF��p��O��^��[0��Bڼ��?\;.x����([���,��X�0� j����y�Η�2CN���/9V!�:|��s}k��e��鏉D(�t#B����
SS��é:R!�\����5 �ZTg*Yт1"c��b��Ѻٓ5z�a�a�w/q.->�ܠ��s����"Ì^���Ke�����S��mTix��j#?F2�Ȩ!�!�����~��[����?�8��e@�������q�y;o�5�r���MB�Ui+3Le���d
�ѱ�̀��g�K`݅��W�d��(����k��r� ���	5H��N0�`�㷤��6+��,�+nA�7��3K�#��0 ����f���6J��%ß���2f�8�v�#czwI�9-i0��I�jy�	B;(H�=r�7�GٰBz����+�a�!�̆��)�ŧmF����+�7��F�	�v6Y���Nެ������,:���RF2��U]y�Ft7Z%��<;��,�q�Sfe�,�,�o%s�@�߳p,�Vo�\l'%6	�岎�����F����Q��i���ĿU`��av1���;�����O��
y��?#,LH\n�M�@H(��R��9�yRm��!c�3�6�� ���W�6�w�ϊb�������8O�� )�,����G�~f���Y�[_2k��V9y9K�N#쫎Q��,�)!�Fy�`�@�J=����6�����,�Bz���-�?����������
 3֖��g2���6�!��)YJ,p��r(��(���D�Ʈ�n�l�y�/}��d �~/q�����)�e�h�h���Xy0x� k�6�!T�+�Qs5��0akR��g�s��/m&ܠq�����@��>@�f�H�����*��P �W�����k6��B@�&dƉ!l�M����,Sa�<�@��U��hNeVr,%6�N��� ��g�q'<��2�Y���t��6��pP�4{��,��c�ɏ��hnu�:��߷Ç��7�츅�"8���� �*�PH���xD���WI��t��N�Cq�E�ɧ.�<$${��.ڕ$%�&��>�cP	t����}�R0�뭥����Ugw��b�`Y*���@�%��"2�_�)���y��f�ګ��.Ҋe�6��mw��r�NPg,M�?Q:�})�7�n]��z n|�x�ܮ>�c�����U/B��v�ԛ��b��R�-������Z42��_2�C �0���9v�k�&���� E��
�"��=�5��(��L^���b�q1�㣛"e��1A?�gH��ǝ�ně����lsw��}�:g);Y�OrI�kp����$۔j�d�� y�7=4�Y���c���@ �9j��+O�G.n�'}�O!�������^����_�C1x�e*A��"YgE͍�J���_/��F�=tC7�C`��.�� �f�BW->�]ؓ�
"���J�dDB���|Ē"w��]�r,s������/����?#NU�^O��H$�щ~���Fa��7�8�)�n�pK�c��U9��Fj(�g!�6Y�% �bږ�d��ы���m���NV��wΚ-Vϣ�:�O����Al��qg��%�^45�S�@���4y�~@��Bt&�d,7�@�1�ꢅ#3o������L#͚&����z%��2�|��<�V邅`MZI>���j�z�b��������ؾ��R��]��%+��rߛ�n>R[�%���뽂<��W�d ����(FQ�4�>��_Ji���A*T���Z���)��v�#�&l���^���Dzqq�]'���j��Gq�$�b����e��5qjO��sDJ�=y�D�oF !:8�{��|�4Ɂ)t��X��)(и Bs� ������5�<�������x9�5�Hh�l���R�f�����-[��.� ��o���ܝ4����Dw��D�Q �ٝW��8��wV*����^y%��w��#��� fe��:�(ϝ�E�$���.�<cr�s$d��i9C�Ӆ@���kw�,Sَ���6� +�=B�B��0��&�51)	����J���멯�b�Yse���%�(8�d�#��P�j�\�=��������"ӝj��9�h%��)�d�H��}U�Q�25Ji�7A�%��|���UF�-�%*c̮�kE��ZagZ�t�udS7�9��dc�4��[��v��"��f�@�uv0�D��v骼����"�ǧ#��[?��]+gS}��lk��]���#���-��-u	!�U��KܬC'��&��DP'��3��#���{�g��$�P�L���w¦V�V��Y=�t�Χ���1�9�	��m�D,�(���T��p
_�E����fy����8����z�{?�J�3�3g��5�L���0��T��"�a���Y^��5J��ޚL�yZx�(�����'&��/uPhc���C�W�ǯ��m�d��"�AW��.,`y.�,̜�Z��|�T2�0�
z��['(����ɕ&TP��N� ou����M]i���w~�:�;�B*6�Y�s~CU�|�zy�{�!�&��Zw[`1�nd���7>U��hK��dž0���ޥѱ�5�� Ɉ��K`xNա.g�D�
�cl����6U�=v�&�C�ř��ۤ�s��I�Q{*U�ߌ
2�ϙ\�&%W^���U�uڽdB�U���l���lO�a���N<��̫�l�FL�ڼ��5xZ���ם��^�~������W��a��U�M���y���f�p~jn����(��g��R�(����3��d�
��Ζ{;�],*�Wm��l���{$�\`�E~��<Y�<,a����ׄ=�oI�=~VMH�hA�:sn�~�{��G�{��٦v]��p2�9V�ht�Mu�!?�Q��J��w1�&��j��#3�t���T��uW7!�^ё�U�l�/�D_�c��[�W����SR�
ڲ� �ǥ�.��"���ܳ8ݹ������<iO�d��ˮ���>��/�.����OR�I"Z��5ի�Y��Z��jP6�xS�?�w{��	�Kҫ@�QD���Ff*FP�8��0�st�?�$�ܡ���9�bvv4������������NJ�h�"�h3���m���5|���R9��t�[f��rO��E������%���"�H���;{����}�L�`�$_0��*[XT�6����b!�ϐ���=�>��E�4�m�Ň�
;
��X�u���VcW�˴�^�/�NVA8K�1��&�i��.FԧV��|t��rUj$���.�f��K�f��a��	��)"Dq��Ρ�0X��bs���V�������Y�w�̪=�Ht����'<֢(+�y�&\�KH4��-@r\��[C);��#4���p�>@��������ҙ�!;ڝ�)��e�?ͷJv���9�l~I6HȮ9�(�A�a42Uؠ��d�7ecm
k�� ����l����Q�eNX��)�Փ=��䵋[��&��*��*՜6pM���޲���oVn�D�=�؟���_�֟�-�"��I��9��8�,���<���̃�o5
3&�%��$���& o�ɗ�'��7�/f�s�v�dp.�Hk���Pw�w@�A��F�~.�4|}!3�?�6��]O3e���*�w�,��ls:2O��<Wֱk�	�xHK�f�:qJJ0_Qu�6��R��G6��4'�Iit�9�ʸ����S��`^^x���>��2�u��-Py�_����(e"��d��b^Z�������b`�:M�K����
��dΒ4���������{{�4F������^���j&�џ{�K����pL�oE��=��z�J2[�B:��.��,4477L�6�p����bs��0J��q�Cc*���J'(̰ec�z,��l!�3�s��9���6�_}�7(&�Q���$�^X��m�YW�ZKV����)��S��(֫Z��l��K�����W\�L"�KZ9Հ�T�~�]�qݠ�[�Ӓ���� �L�$�0#V3�c���e&:�K>`-*�?�:eK��OԜX�`��ސ��v������)	��ε��r����´"��̃��|'�,���|B��p:��y�Ͽ2`ka�VJ��z��(Y@OV~�2->�a��PN�|l3�.� ��\j�P��e�'�<��m#g�s���94����U�ԁ�x�f�v��]р��u��aD}7i�a?���Hq�qZ�-~���叭"�d�މl.�u�,uoC/fV�Z�%��<��X�#����p���u����U��@P���u�	�%�T����(�
`���`a��/�=\a�4�Nb"�,���z�1�'���H�3m��bL�c�ƥ���U��ғ6���+�P��9�j-Ư�z}&q:��R�f7���ϩ�-����;����쪘�ҡe�f��)Ǡ3C�j�+P-뇈�0�U��I�weUX��?Z������\�= $=A@�B�����t�QT�`�JDG�ZFY�#������1��BC��S����dZ,�e�qZ�<��G�q� h�I2����aI%��Qo� xb=���#���ʬxWC�[X��	W��Շ�9��q��B���O����������)�l�lR�͞�K�������x����E�us��\�-��ܫ�$����Ҳ���]���j�G�w�$��ʫ?�*�u��ڧ�6�G	q!X
�d
$0��@�u��M�@n2 �#��V ��֎i���Px{�O	��ԥ
�`�KR�,�<�zw��t��e�F��z  �.ܞ�u��6�D��HʿDf����Sb�u�
���޾�&���t`�O3�s�����ȑ�E�U��bv����}c��> �:&��h���9)����E#�X82hVU��_�H�Xj�=�(sWeݞZ��c�b�AiI���&�+�l�^��Hp� ����B�hC��'��Ә���E�lV"_��{y��7�ړܘA��=��_s�,A0�E׫w� 3�0ƂZe	Ć���s
_7̌z>;b#%H��Hx�_�VG�@r��~w�$}��� %��/T4���q�|u�t3@Jy�w@��<t*O�ԗ(���	�
���D,A�v
�*1V��Sq����+��B�a�pB����$���Ѓ(.������qT�N�U�6ɠi2�-�^���4������U�S����<��hǮ�nw�*��	���}շ�frrq��K��&@��Y�w?�u���>��H��~��@2����SI���(
����rB���O�T��\A] s.��	�}D����������PQ��㲘�c�tm�:1�8O�N2��4�j�*�$�.iD��#��G���s��3I��,�J�x��	���m�4BۉS�G������~��5o�ѕ��R�3�H�.���w�[��X5�+�g���+����(��_�����)g�`������\�̔`0��ĕ�(e<���	'ͤ?��6�\)b�;�hP}g���ˁ3��F�� D��ZM�8�)�t4;���ʸ�ɿ�thJM2��u-�:��q�l���n8�7NM;�S�Dm���cQ�#AX�=p���LYF�u7IlM�]Jf�Kw��ꬦ8��B�6��i�ܣ�ԫkS�*�H	���}N�8�5�K�,��_�"���x:�~_��6u;���*��d޿��N�ʩ����	Md�%�����cV��@���E����,���|t>S��À���^��$i&m��4؏��<Z���e�����˄�e�K2�Bb��rN)��L�jfDc�F��@e�Pe6ۨ�<�j��ȃt9�J��PA��Jyj�[�<О}G"�V*I$��u� �p��V|Xɘ�)��h)�[�����?i���)��VHe!��{���^�	*��q� |-e���%�z�W�w2��4�$$�B�X�J�s�C>�Q�ƼQ <8h�gG����8�=:0�7����,��=b����ow�´�zp%�[$M���˛ ��"��>��VG��������>����jE��5�ʍD�= ����hz5s3���</t&E��@QH5�S^}H`��?{N�^�gPK����r�z�E;6x��rQ.��}�S��䛃�G�8���|o���?��O���m�r�@��f����)�u�VlC��/"7�%չ~���`�����ꦡ�( ��&G���=�B�ڰ��E �V;
�A�	���I.�Du���+·�F
��Q��M�a�`���P��~���?`C�Sq���C����M��2���R!�vC�y�]� �0#ؤ�[�֤� b��b:��%:%��f�p`��}���ޣ�N�]Y1D��2�#zٮ�B��>����ԽT��IKN*ɚ�}�M`�v;��^<�c�YF&B����
<�Q�Pc�d^Zn���P0���rs�����Kđ�����M�/�,4gkoMv��<M�4
��}x>��=po�WS�H���ZƎG�s�_+��]�Q�$9�'�E\�l������K�=3�:y����f���/5��<l^�@�QZ#I赏���M�� �/�3��8)�P���**���>��֥x��ZŝAa��?�Nh�\��\��}e������ƷdZ�G�J�3���fi�W���]��O%�0�,9�'Iun�̩%c.�t��L���M1�t��OD�19Y���ϊ�\�߷�	����!M�<]K�?�v�pY�5Mq.����=�x(�J1/?�i�j	T�^����gK�!X�@M:ro�V�(�y�߹��t��D	�r�-s�S��)��<�g:�;��0���Y��n�Z3�D J�V]���t U�C��F=�"�z.�[IEf��^���j"�&�mX���t��T��t�p>]^��0�o^�,�:	�y��+Q:�"���u�'�A�]���8j��^	H���8�OX>�b���?���#p����^L�44M����d�$��^G*!��
� ��@S�,�kZ��-ޓ�g �����4�����:�����[�v����f�Q\ 1F�,�[�:*>�=�b�qV���#�N��MU���i��_�2!<v��7�] Ý�m���%�{�/�o���}��H[����7��{�ŷ�7�66�Mf�mI6P�7L�Ji
,����(8��{1%��S���P����Mk���N}1�Q��w,*�,�O���_��l߀KM읥)9]�'0"��T;�6�Kq�R�ݠ�xR�_�5xdn,�
�S���|P�N���������|V���lգN��b�ԐVΕ{�L�c�[�ćdٯ�ڔ�3��F/�BQ����:l�P�n�J��C����$����W����r���sP��do�E��Z���W����/?�:����=�����Ŋ���_����1�-W{0hx9��y�,�0�򏦸Y���'-:x	���08&LfXc\p�����#hh���:46�ON֯n���<e���9�,G1$8�ۜb����Ͷ�C�8̸-%��B-�dz�M�@�jCJ�J��tG{v�i�%��q�y�'���q��2����@�@�v%M,��Bw���km0�,��4�*ԫ��z'����.��-,O����e�G�]0��cw��ټ4��M�:Yz\W���
�m�;4[�~
���ޠ~K*|�a;6��Mϑc=q���`�u3�=�R�2ZmP�ևJ:�.j�Ux8$B��e�[<2*&�-���ǯ߯WH�ac�U8%\�:�5�ꓦ,R�C�J��5;��F ��C�	��&Y�[		� ��u`�/_���6��Ψ	S�X�ų�%kpM@�1����k��}Ú_�$po�q�J�O�bL'l��X`�vLd��9��s�Ofr1W�3�Ij�d�{�g����y�=����L�98�x�	¤���d��*zm��A�Լw�	sת�����5}���|-��ܫ8���VTb�8�ҭ��f$I�!K_�Lj�׀p��Q���_�H2�۾���E�v��&�4�i����f�N�v��y\x��/� F3=|քy��{�NRnr�'��R���n����x� �78/a�(�;�:GU�ƕ_�bQ�z�V�G�Yi�H�Q�	n�a���ք_@�?W"\
\�Il��N a��|n{*~f�_J?��
����M�,���;�r�l����ys�V�{Z6 Ś	fSV� �W3;�亽�[2��呲�������*�7�� �������b��l54Ԃ�#!�����N���&~��	��X�NOK%��3�͐�~��Z�@�?�]�l4�{���*�`�����*m�X�u�躱g�u���rW��6f�a2ɨ/��և��$O}1�#�j��q�5�9�V(5����E2Y)���o�ɵټE6u���)����PG��&�`{%�B)��߀��8�k�T���md)0(��G�]�9��,r�e��V������v��g�& ���#ڤi���X�`�� �k$��aM�.B�ӷ���H�Oy�:�1�Z�]�hM��\�?��d����A&��Ni�Yâ��ͩ!ND;���*�SV�0r̥��W�$��e�؜���H~(Ɇ\cx��d���4ѽ�3PQ�ڳ��z{�..�/���Q�]�����r�G�/��e�����#6:jb�X�Of�4�E�W�(w�f|S���󗽬�U�u��y�s��A�z����5(1�=�N��a��"x��Q�t�J'Ѓ�p�g�'HB��p��)��E�G��Ս���F����9h�V���v�cX47����g��Ի�
��A'��P�.��g��Ͱ�.�WC
���M���"D�B�P0yْB�x��'�H��"��,l��;^Fux]�naA"j�oT�ـ8�!�u	t���b�ψaM	�	�0�y�e�X���L�í�#2�}r9�
��dw��8�ۓ7�_�9�s��P��6��o�{?�1�+����W���6��5��![�I���m8�@U�Qئ�+酞�H;�q�$�tP��JP�xY|�/o|�e�h}f�!�2�Ή����XK�������C2}�%�����ܗP]�x��r�1ى�R~sC�� YT�) 9���[ax�R��l�7�Q;������5Q9
�f#�<*��N�� �t�0���.а���9�g݆��=��˒�Ԏ-�դx.)�_�Df�g����T%�"�>�ڴ�3��u�����>�a�˃�
Rb���N9ԡ
�}:kˌnK�����;��͔$/���݋u�Ӝ��͌�
��Z$O'R���ڞ� ��d�ѕ��Ocu�����Y-����l�~$�8��HS^�i���p ̎��)[I�y7��B/~�~��'v��Hq2�M�A;ݼh^�����}&�W���(�(��\���S�$�,��V�(��y����!��x�0H�E.������4v��s-]��rj(�D�+�D�sXf��H�r}������_��m=�Ij�OY-�$)�@�]����/��@�pɈC��}��{.%��`D)9VJ���F���&���iA"�y#z��]�B��s��YN��fkwD�m�Y ���A�j���*�-�r�V)��31��PQ�̲�~tN�3�u�X�)E�W���s��]���Wj�j�:F��{o@�ȍ>0�$��Xm��&� ��C�F&�}��
jz��6�3�0�~Y_9R��H�20�!�٥�d����x\���:����b���F��V��;-l� �)Q�T}��FU��V0�_��S�o�zݼ�,�]���,��i�՜����NdX��:�)g`%�@y��`%0��?u�㶈�g�*W秧+@U4F0�z"�b�s�A�b�%WJ ͧ[�-J��)����0�N�[Do>��Z%�U���ifuB�Y��*�����d���EK��R�
]j�et��N��
B�gZwt�|�-���&{e����k%ԧB�b��p/vq��޽ \Sa�`�#��f�g)k6B�����-\�9M�`��O���$5���o�:�dzʿ]9�U��
���Jv���5��awP縋zБ�V�Ɖ�ְ�8Ә�_�(�+n����w�*�2,�U�������W�KW�⓹�}J��а�G�+{U�S�^��6�֍c�I/z�	=BK�_{�.Ճ�r�/ġ;��|��ؾqD��26� 7�҃��jو���ˢ�T}\-�a֛�mfG��X#uO6�N�E����*��{����r�+�nˡE�bH�������f�g�H~��(���oS��e��R u���"�z�0��&��z.���Ќ�̢V���x~칖��҂�_�Uo���<��6`�X�R��R��w��-"BD�Zm@��-K4����DkC6�}�:\�BqN�]7�v6��]($�r����2/ɀ�t�u^�W�-]�F�Ʌ%���b�ӕ/RX��@�!(�X�&oR��Q9�+l �����Y˫�M�46��̼Nx�		����lP>�?1+w'^[@�b�1Mh*՟Lr��V�͛Xp��Tg��i<.F�+Fl�&G��/�����	d%�U�����{7�P	�d
��k\첅�M�6����6aE�ahOV�F�?
�X�(�m�_*"s�9�Q����J�Y c�O6Ym�����	����k���2�ye_7�;��I�5q���햇�6��1���(���]�˜K*{#qP��g���7<���̨��mM_�in�TS�k�����i!l�ia�����N7k�=Ę��0��~޿
uC�~����ʶ9\��S�+���=���_ �y%[Aa�D��3���,���jdb(�6��f�K�<F��V`�Rr@i{����.	s;�ΖRq�	U�HX���	�����W,�z�$�ƼGT�QS;�h�kd��� ��j�j񇒴U�UT>�V�q����;�K��j��Ӂ-<�)A����r��8��Nɧn�Q'R:g��޷�9�L!9\�_�8t�������l[PA��ߙW���m�#3i��������JZM�z�ȝ�Ƨ�ۆ�d-T`���J̀��Q��nٜ�Fk�luC�4x�i���^�k��bp��;�V^0y�W�� �0@�%����S4��/4c��{W#s'=��jఅ�;�]ˁIJd�\�n	8Yƞ��y%G�-�O�{��!89��aλ�1�xr�謨����%~��Uӵ�yK��]�J�OS�Wl��Ւ��yD�* I�S�vfǂ�<3vqNx��s:�t$'d��wyF�9�06�g�;��jLd�{�_"ݱ��ޏ ���r��C]M�J����J!�,݊�k{�aQ-湪��2+���"�R ���-��]��^��Ɓ֪�ko��o��l�v�c� �.�h���PX����\V6�W�)�l;� �����=���U�ւW�l18gw�c$�4`��<ַ_�{��0��=������}�s��%A�f��˷R^>?=�uK���I:-��R����z����W�id��t(���L�uTbI)cʓ�F&�0Lx�5
�� �
)W�<��|h����s	X�t�c(���R;W��m�-!^��80�$1[�?������<g�!ȼ�%�����/(B6�L�'N���H�:h�]7��3Y�^CHc<Ӷ��pB���/Z>�0�8�3�����1R�[�>?��)�

dޅ�/�:@��y�_�����'��)(�����bI�w��e�J��W�0�m����:G��r���u�9�z����o�uH쌌���N2 _ŘWJS	���8��^��˯T{�gKI��E�����t�q¢5�*��G����P9��Du�tٙ��s��=��dr�U�bo���Q�I���J�Kt�&��J�Wb s4��� �ʪ��.�ow-+��|Ȏ���f�bD0����*%c��3�w�/�V�>.�ku�8[��V<��� ����g�r��J�}�k�'�8Q�s#���k������8�{μ�̖��\���
�� �Ixu'5]�N��`T�FnrGe$=7�Rڇ�.1�o�����;���{��*�z0��蔃��a��/&���Ϟ�۱ᇲ�E%B�_)\��9g��L�A}َ�� �B��f�b�QE�F��gh�M�b`���
Y�p�+�h�C;j���\�s;�s}`�4���'e��\��tc�xA�AFr��xr$��Kc����|q�Q����)�-ՙf�yp�Z���6М �T�;ѽ���z{u�cs�ˑbJJ���n�V�>}�vӂ��`�x�f����ңU��jo�p"e*�\g��P���'(l��i��֮��W�ݽ���ڞm�ш!5����F��y�{Db��i��S�u`�lI�6f�	X����8�͢��Q �>^�g"���!>T����F83��!BA��˺�km��/��<�tBw��s>O־�e� �몲j���?Ec���^z�_VN�0��0�l&r�GD2�<j�:�,4@x�gbX����E[ZD�_��\�φL���0m��=4hlb�⣳�5|&Jk�#�
�����}x��,�N��6E�![��2#�?w���I���Nu�H�fGHf������y���m�1�^�ձ���HN�m�M .C��u�/�0(�j���JpD�!�)�Z��WHA��*���jǗ U���3}$^���D�h;&7G�p��"X�#vk��xQ��$�H�N���!�;�a4��H%�B��(��	G�z�R�:�3�8�#�0yt�*��C�95�9Rg��H�����*Ʉ�� �����E���*w�����P�Z+<���X$k#.��LJv��<�������ut�����Om�me 5��Jĵ��#A�/���FCठ���:c�G�g�
ΚD���UP�e��du��ٱ,<�-j��2���&�4�6�CC<���u!���r7��I�YeCc�^�ܭb�#���t�I���2�~<��~�� qJ�<$t���BM���8�-���s�eF��ց#{h�!~�	�й+�c�k�S?H;�V˦�[U�\ ��<�!��md0e��lo�1pj�f||W4,x%��n,_`w����qv�H���[fRn�9����loo���M��E�,�w�|���g"���k�#ڱ��1���cV��Mt��,��l1�Kxa���gO�	���=L���~��Df��t�2�~�P���]7NJ?2vH&��� x6���z�=�v�m*�D��R2�@5|G�Lh��_�	<CL8�29�_k��H���k�6�>�DI��PC��D4E��/��	���~��s�n@xY�o1�-�P������ބ���v~�ި� �Tx����p1��إ�J�W��z��F�@��N{�)a%/*�W�Q;�[�M��+�{�r�[� -yF������4N�;���m tL��|��Z��;�гD/_����y���AD$u�{� ��)ݳY�~_U.�#�ԈT[�ʗ,h�a��	���dG�, W*�
_��`�f��CGDL����
�bB$��::g�Ǡ�����r"W�FEc|2BO��HK�jv�p��9��[˷0�tq2���@�gEV(Q:޸��Ě��7Fv8�(<*w��3��jgF�'��n�!(Ʉ�EK�h���YpR%x�)Z��U:� &����zrR�Rש�A>����I�ظ�<����`���<�H|$�����"���Ân)Tܶ'�+E,��K-�'��ױ��z����0��}N[����P[fc��Vm��&(y��׀=8�����/���`E�y������[��Q��(i��G%g�i�Ƽ:���+�o,Aм�Zlj�@�ob#�vg���S�s�#)Z�Y��L)t�a�Pu�8����-�u�b��B�%|W�'��d4��H��.�2-G�w`�"ؑ�w�����j8���nʤ��0�M�0�<�+� -��<,����uP�,�c78�F�����~+���)�����.�W�G�0|��QZ�6�=e���y*�d5�Η�_�H㻼Dn&)��}��&��WĀ�F!�����$}�9W����Y!x�~?�Օ��I�vb_e�ֶ�CE�i	�8���K]��~wcn�@�$�u�"^��o'B�\GC�]�h�.�]B�"I�P�O�D�|��b��4�C�+����s=�mgY��P���զ����/�A� ?�?�8ǉÓ��	���3�rV)����y`��� �]���X
,jU�����_��op�N�BS�p�x�}����\Y��+��A0�Fl�" LZ��^KA��W�ݪqu֞T%�,�y�y*(�q;�l������>߷����K��_�N����6������;/e���t`�Y&{jـY>�M��IGV$2����I��#���đ�AT���G̽J����
��#��t�Rsf�Q(VH+�Z(��4�-{@�4�'y��c��4��ʎRᓡ��v����̺���"���F��6W�E�-܎��@c#�Ύ-�]bG����p���rc�����Yv��v��o���^Ņb{0m�L)�]3�d_�R�ȹ�,����>瓞4��;S�_]���@R�����[�����ߌE�Џ����jq�Wt�/h@�X�XR4���Eߦh��=wUluFŞ�[p6�?��>s`؈@r��`~ʣ'��7�tP=ί��.S�.*��D���f��Z�&?��j@��.��o��#n3��+!�-��ʱ"�X����GWe��)��`U8��Kͅ���4�J��79[Ѧ� |d�:�����s|l���Ka	Z�Fk^?jPEr�4Ał��Jw�q���\�o�Gs]k"z2⋮���)�a�s<9֥�.T{�뼲-CX!W�!-'>M��KP�C1�
%��P�I�ʹڊG�	��v/���^�s��a������X]��6x����L�2I��Ȇ��"�O
-3�re�SGu� 7!̕+�f���*�Y�Ć��b�Е�[�4P	 �J+w������u{���bH�]���u�0)�8���5��7	S<f�#��b�Z7вZkb�^���
=��1<�{�����B��q2Sa
�R1�Z���`�U��zey��e����sȷ�:f�4�;�aRw��uVW�`�p&O���U�����"���w:���@2�LV���'�a�n���:E�<�GR�g�������.]�n�����[Z���	P�`�Z!�	_�^\"so~0x���0�u�+�E��Y˅r����C������݁l+v	��?�guf9�I���fN����XH�Oq� �0��;D߄�~d���3p�VI{G�(�gA`���\�zY��ۯ���]b<����eh�*y���aN|+}���(�ۍ�b�$�zVb�g!����L@|s0�4�\L�'��UY(��F?Y���5�|q ݷ2�H��<�5"�SFȜ �@΀aJbUN`���Hn���H.��f��z'����}�Q�����w{uz�Sӆ@=���e��j�Q��;> x��$��<����P�1f�'�n�`�Ų<�9���UL��sl�2�I��$�i(<\��fL��z�Ke�M���'ȟV����˜����nN>�f,��q�`;򣎒�7!�׵�W.c��*}}ȍ��PoX.+M�/0[�k�{����P;=uz�S�x.���'ˉ�s��~�=}����U�-��,�a}���* ���ߒ��܍�Q���kV�Ψ�U�}"Nr�:����qVwt�;�<媷��Q��y~��J�n�2B��F_�Q �P���3Z�]8�1�sQvF�oVQ�÷�km��-Ŵ���P{�
wެΡ��S�.�%��C-��N����.<(��q��}��t/�ی�8�Wc�n�7�#�KQĪ3X�&z�P�[�x�mVС��b%�c֏���&��q�����:�oX���8�Z�W�s���(Wb�+�bѫ�TJ��ܠ�ţ�6[FJ�kzBnH�%k�&��_zm&�����YX[���Y�sr��)�׊;��I��.�V���w�.,�6�aLT�}�r���͍o�� ��w9��/��ToJ�H�v��Q�(~�`�3Rr_���u�2La��4��~O��А9�ԐB.7���|���O�3:�ͫ��$B2�H����8�l���Ȥ=W��i�Jzz-�?��{��]�����[kqR��c"������	��]�55�`xZo���I�u����s&�{��e9Z���[�o]�3���r�)�b}y�r�X�c�9n�lzj� �"F��3��S�x���.�^_G(���x@���`�R`��$�(��h��J�Є|p;�H�e���&Q�xW���;�m �KmpI4�9��y1����Cepw��*��A\4���l\�ն�#>��̢�x+�k��dЩ�Qq�*dp�v�K�o�ܥi�%
�8�}���^����Z��/�!\Ls	`U*������	s�g�6ԑ�q>hGk3�b���M��;��ʈS,	mnF�;"��p-�g�"sz�9�.V��W���s�RrL N�p�+��� ��X�0�El
K����/;���AG��Z�@[�D�A,�M;���`�O��k�ң��B�m�,��t7���W}��h�"��PZal���h+��X�b������p4|�@69�1�	�X��_�4��W7��O�����L����*�.~+�>����h۳��r��]�K3��N�jXYE�����h}{��C6or��a �nw�Kbi�έ�m�������?N��(�X ��F�� 0�旤k��	A/�WD�P�A�-\�$�w ��JZPۣ�_ݵ����PY���g�?����#��"�%$���H�~0D�MPD��健~�������y���=n���T��+a��ޡ�y7T{+*����7�bG���]��6�������:�(��%��D��!�;�����T��y��?- c�Ɛ���+��"a��l&	����p�E��0[���dV���TSֱ�or����g;�Nk/E!��` "pW]��n�B���T����{_��P�'Yp]�e�_s�
�I��9���Gi-x֎��ta�`�j�"AK��O�:����:���mb���B�5�GS�Aְ;:)����I�Z:NǕ*�;���!~(4	4I�y���^~�_��/"u؍�AN�� ʚ����.�|��'�v5Mo�	�_p����,��~*+�7W�ŗ�  &�M �� �gF��k扭pfkǙz �Cy[Xh_te��	����
l@&	��#�֤���f�d��^@D	�i|�z��i�뵩m�(X5�x� N�12 ��B~m�2�mpl{��Y�
*$�Љ(�&	�Ik/<�� �\��n���]K~�4z�5��N�ky�Sғ�� 秧Y�עQ`_b/M�;G�~�r�Ne���;��3���r@�44�U3���mu����)���C� au���ыt��w�$ߘ�Q���`_�:�	>%R��S]��M���\����u�G=��EV�.��X�Q���'dM{#R��7SJw>�3t���㢨T[�$	K;�b�]�E�\�|3����I������OI�L �]�q�M�A ���N���[��'���z� 0�~���*�f�x|g>r��Ek -bא���,X�AL#�ª3I�d����[���T/�5�+n�����ӂKyG��U����Y���IT�Vva-RC\@Ao(\qv&�B���I� v��4A@g�
�Rp�>�x=�w>�neCSU?5�M�_��E��X, ���1��;�xYT oҀ��L�_���n����%pq@i��HhjR�N l5oS�x�d�W3ő��:��8D�����PX�8x[EO�h��y��D^'am�E����	�ݠ�"!��C�����OB�&���,���|��ύ�^J�����s�x0�ɤF��|lN*��+�F_��cH͈j� 5�+n��q����|S���˼	��d䆳�JMh ��lFN�ש9TlB{�	{Ƙu=���#JhQ�FT�PU�FN?cYߟ�Y��"+���4�m18}lK����2�������]v��aV4@��aYg�i�v\�To���聣T����x���l�^��
7�u�m���.�z�%��!�|����-[W=�är�dUCp�d�YJ�����/B��4�[�.�}Ng|��o�
��Т~�����N2��72O���ؐ|�T�%$�:�^�Y���%����[R���O{�B�[��Z�Zm�@���鼃�1��u\+�/�]5�i`����P�;��,jaq��<1������eT���?1c����V�W߶���˅[F�K��Gf���t�g��������J�~F.�B�'[�"�bƌ�BA;�=�{�Uy]�Y%����F=�}^��5�-�0�>ͣ��Bm��P�K+.���j��z�=����h��R�3�6��bK| hj<NE���mV�	c�*>���ѿ��/a�׸��jք�}�?�|���-Q���iבl�����XeƄ:��L��24uW���O�_�Ѹ�Sm9m1�֐0�z
�
������$�X͝B�%������v�P�<(� �I}n.ͨa|����< ��l���.�`*�v�IN��0E��k�q��ס�*0��'m����|�x�����N�pƠ��)�2c�$��S@6��*�+T�*��*��z�XW| &\x�|8H��X����y?-����n�{��HZ4wL�l>L-U�w:'m�ɔZҳ��}����Q|��6�s~��`*��
dYz�N��+���
'�_�p��Z�C��s���`�Z���TJ����`O:S�L�Α�:��Y�Ģ)q� �X���$���.0�X�C|1��%�����e�Of��=�C�@���}9�E����XC �����b�-|y0Ar L���g�|Y����ҕ����zhw��9�j�8���(��2�����Uk�,�D9Cv'D��K��C4����L~�
�^:_��w��S�ڸ��������:��(��HV&x�k�Qp��@	�81d��}mO���7!&��xE|{���y��O��}I�ݧBϊ_XZºळ�#)�ͭy��Ff�໫�;�˷ZS��Ӛ1�{$�E�w�c�nt�V�~�R6tܯ�Q���j�ΉF���_6����ɒ-*�I瘹�򷓔���oUb�Y��N6&$�a�ZK�CDs%~�灉�7l@#��>��%ds�b_�ެ�L0Flm�?��N�l�,�m�*	�>��a[�=�S_1�9�/�VI��Je��T�D{U.t������ a��&���0�F�X�`{\(6��4����M?�����'�`�b��:NP�JB��ʫ�#��q�_r#IW�=�������pxW�
�ܫ;j�H��3�P�ȇ�Q�8�L�v5�0C���b0�T"��m�ØG"�(�Y��{��ɒ��;dL	J����$�Z�@ɾ@��ٝD�s���P���"�'kD�x�*t|r�O���P5����K�՚c"�Y~�>�2W����&I����ɷ\n�N�,X��Y;>Aǈ��!w-���4�x,�����ڙ��$��ͧ��z����9���է�]�((�H�~� +C�h}s\��=��&{(H������#�>��6�A�ŏ@�H����Z~��b��af��$%!�$m���-�h��$|	{\�N��1�����Ƣ)�����G��ri\-�s�R���^
��*k6�r!�>_��n@�L!�����E�>m�]D�A����!�zy �N5v����Sf��.�������J�<|-�x����I<]��7ސ�,
�F��(�i�[�Ǿ��M�c{�6���&(Zfʯ���2O|�6DnS�{�g�h���Uַ����v�1 A��p���(0� 2~HZ������Z�dfl�x��T�ʢbE|9�H���2��aΐD���"��L�+�	�M�l�3�a?�>����$�&��ؒ�TH{V��Mz�:�숓N���� �-������O�#��]�G������@���u�0�,��q&֛\����t)��#�5R`�g�=%���oa}~��ǃ���,�ҩ���qj�_ ���)���}�'I�ʬmo���,���ń���$����u�ӥ�+ 4Q����i%�a���8
 {�d"�t���`��8&zeΏ.ِ`�q�Y<�J5�"�mI X�3	���9}#Ҫe�����Ȇ�S�S��S���H����`�
!6i،��y�6�ItL��)�r[����p��I4nm�pƣ�.1�*�l%6' �)�fؐcb�n��-�74AMU�����sIݐ����\�y�-a*$E*斏}�J��T�~��B��Q��/B �,_�"�NTm�b��?|�?�$)�S
����ۄS}!n"���Ĵ9����t��.�s������[��į��@y�����9�Qe���Ɛ�?�%�CE�R&��'BY_g_#H�"`��&&�d߱L�K�H<�vDK��X-��1����.od���$teؕ�HN��.�{c�bT�V� v�z�;*���S�Ǡ:I4���6�����U��&�!��Y���	�ϖ�D i�h��ӄ���F����rm��� �WWs���H�.�b���}->�^�%�D�hY��/$(W[���,葱��)���������t�{�0�c��ٝ^x%�j[�{�\�o�)���7B�ĳ��ӳ�_������+7���:Zu�)�jh������Y�텔��l����
A��'.1���K�b!)9&� ʗ�5�X������:����4-�ʦHG׃G{aϑa�d�������ϯ�c@O��;��zb��K�0��%��)46�	�p�LJ�)��J��m��h4F���(�]#��8��N�z����0��j��1�n��G^s��[T.sX�C��q��º���/��Z�q4����-@�쳊!������o������L�Hb�2c�vTL�o��˭A����#������D����!�V}Vj����T��K~Ir_@-�L�ׯp���y�L�s|��,��r��^�9G�d=�9\Y~��]�LF�,B	C�]����{��Sa�H�%�+9���,��f&1�L�]ǅ���8>!. �%�"Ѓ��8V��(l��#�.ɒ��l�3���:�a*�=�8;���]��@?�ʍѾcx�[i�e	��)�����y��`�q��t���ߟKv��bX���"�X�<H�*YxщM���cp$�|��eTtٚ<�{��g����� Ѱ�Q���:�%^����uJ���D���4:�<bC {"��0a��|�swׄ���	������ ��/u��X�[:`�C����y�P�Tr.}쒩̘.R�:� �o�� �J�[t�1�_v�rf��|�i�q{�]��_�ˀ�b�$���S���7�I$��J�$�lM������Q�Z��x��m�5G�կu0���g�!X����Mt��S^�^_�m��j���'ԝ�������b_U������P��� .��e ��+��	ǟ1�嵛�Lb,�Wh�
�VҦCK��#E8uJ�"ߧb���V�o0s�z���?H�ѵ�}T��l�َb�M�.��·T�2b�q����@	;�3:�3�i�!$�c�6ݩ98����Ƈ,���P�Ys����&�����$��m�{�4� Rܮ]a���?���r�Qt�_[�b�d���C��\b���0��i�����F�����w?��:���H7�Bv�ǖ{������j�V�J�#�Ց+�\^N���Y���7x�C��f��Q WB��F�����������8!���k��.�9�q�SY�h�~�e^>Y�Ho&�ԃ��j� 6>nbw�`a���0q/Q�̸
��2�sew�����w�.�x�_
�A�}Ľ,ߕ(t�JoW�Q�y�eN��a�"3�������7X���)A�+��S�=�&dS!>�!�׊_�M���)	�2eۅ4�&@	�� �ޞ!��/q����"�XV��e=Z���e�Ԩ����;|��1Ύ��eܾ������	Fe�Q�X� ƘTe��u ���t7�De��fT -������KR������>��Ct4_f�\�o�|��*��sbp|�����E�"�o��6�_R�k��Ml׆ MS��s�P�� s4����[�4Vl��� ��v�RL�:ݼ'��ga�&H��w��V�㼡��m���h4M�њ�y��AnVJ�}$�GM�)�9��5�?������N�V�%�NB������ 7q󋮻���T����O�q����]�I�#|��I�4������f+��uf�`00��"�q((|K����T���ڪ҇��`���i�����r�Cz�+���*�4�M����z+��E�;咥χRِTy�(�f&��-FLStC���|ťW���I#��n���4��L+Fɕp�\��t�"��*.<[{R�U�������߀�_��0�]��[�8��5j&���#�_u����)/M�},��<T��q�.�q{4���,\lU�Se���
z�=���z$�L�Yt����z�w
o5=z]$ x�g5һ�9S(����Μ�2�#�ɔvv��Me�,\Z�z��}+N�������X�oex�3#U�����Ɗ_v���n����8��Y�81����[�����xѱb�2�.�v-z|KAMg�C�S�8�d |��&����[��#Y�u�m! ��ǟ`_��#�'h������'@]��0��A�;R���Հ��^� �j�z����������ωp�n�

urY��Ù��m����_�-�=�����]��.�7�i�J�$�`F��'0��^ھq;���3��l������u�T8R�*�EnK�zN��K�ݻ�6�(e.�S.�����7�Eڮ�X�9[����\�i���tDrO�j�EŖHn�����r�	�M ��&�l fp���׍\�c��Q�^Y�ٳ��ĵk,n�wt�B*�2��@݉#��%b�-<ٜ�c�3I_�DM�7��&pK�����8��E�r���D�U����w�Pf�H��~>��S6ɚAtU3�_��y�������#2�����B-�zz�
��D�(����(�@zѥ!�������P3�k�9f�eOP�z�#}�=-��ꪾІ�nm�)��IȜ� H�U
�\j���	}���q�Q�$o��������^�j%W����/$G_Ds/W�x�8�Ff��}]�j��a�4�t��t`�� �F�P4�ͱe�IIx<��	���0�g�QH�����J�'{��(r�%�����E�"Q�[s9� wc0F�$YY\�I2SLQ�֐�AY���o���ti��W ���]7i��n����� [�|l���5�+�O5�%��`�|�N�K��RR�1�/��mۣ<I����L�`���-5���,~h��ln����`�۸�<��o��^t{�k&�d�>�=D�nP��
�z�����g�XϢ7��i]�{�D�oD��{� K֝���ؚWY�	t��#N΋ɬeC���k픥�.i��g�j-��fڹZ[�1j�%0٥&��1�6���e)��ߟ�q��q�[���k� �D0�G�L��Y�|ʨ�S���WM�a�ַ"�� Aw�<[k;�Қ�@�	�R�T5�5�ֳ>\��j�;�W'	ːh�.��'�k�poH��.��'cY�9�`H�i��|��\ClT����x�i��Pͦ�K O9z�\�!C*J��d�����,��t��J�m����[��{���{9	��G���p������rڗ����%<Crކ�jCw�c��=E5kp������[�$�\�T��EL[�K��I�"}'�>8�A7��<L�J����1O/a��M��7���j�	*_�IG6��TA>H�G��2��铊F*��`�*�rT��h1#mk�����\��P)�/�/���_�3b��(�X��k��]��H�B�Zi�����l#�)��w/�m9��>�5�����k�F�S��
�,����
�6.�)\"H�f�ٱGB-�S\�{aa�OW�>����U=6F�E���dؗ`�d�k;%g2����IR�I����&]�W|�Zg�ƒ�K��aǖ�nuk�'I�����W"�������,��6�KL�i��i����7��#
������M z�����M/�	�;#_�_�A����Re	nF3Y
�}���'�{o� Z�[��5��W ���$cR�h�Hv�%�ջ���a��iL�cŴ��J�[�J�Ѷ��m�5~E��]��6]h*�Ŵ�0J��(�%���oY#Gr `Dl�n�,,��\�)�t���X�D�F�E�.f6\l���][J���W�����)h�`ޚ㦒�%|恕U��&�m[�{"��B��-�8O��n�֐;��x0�,!��;-��W��p�F����mKd��	̫t��n���T���4�+^p�FZ'����}+��4[�~�SMY+�����r��JY�y��>R$)��J��L(��
P:}������a�9Y�:Cmf���Z��9��������P��<n��&�t"�8ҧ��k�/����W����Q�K��}��fO1�ǝ �U�<t�J�",B�	rVg?�m���L�X@ �V���� �s�����Գ�DτZ��������;���$꽺.=��iC���0�|� h�4@xt2I��I)��!!;�*WW/��`��G{���CƋ�w;/QΣXw��&v�R&s�ry0�x8��SY��l6�/\<���hK��{�ԋ�M!�F+��2	�&�F��V�ynZㅉ�{���
}[��+�dI�~���Ȱ�]	����3��;J>��Ô	ĳ9�𷄡�J�3�[w��!ߐMk`>�6���_ئ6��υ ���Q�����^e��:�N,B��� ���cwX�ha$(Z���\]��}�EҌ�K�.�$Ê���}��FԲ#���Vn�c� R�~4[m�)>�"W>]��B�"�^N�2�C�(��n��RJu�	=v� t'&��>�=
���~�Y\4�! ��#��%j�aU�h���a��C���^@3k �/DGl�4���X[����s�.�*����~��</���l�Z�� �?N+'4���q~����(���'��\x�*�(���	:#D�i�,�<�ߕ#~6e񐌩Ko2������r�+�r/��ʓ�|z��l����9�Y۱�uJb���P?PV�j2�;��;�5\T϶�A���uP!aM��X#�����4TqìcE��,����@!eb&� LDP���3E��,7Bx��q
u���B���a�QS�pG�u��ul;�͖��Ӡ�I.v=^sc�W��AbӃD�qe!�z 9o���E��rפ�Ҏ��.Α�!�Π݈�k�]�{��:�:������,�a�D�I�C�9�����V
�g�����f}�������u�Q�[��9 �:����E&3��K�Nl�sM^;�<ڊ��bb<N�pL��%��ߛm���o2�Sְ��X{ؐGu�T��yB-HgN_0��lţ�M�y�!�a�/�I$�a�~ Mٕ~�rqs���n�*�5q2O$��}��J��	#�;.l��d]��ٌHUMJC ��������4*�\�@�*-�A����A4l�HZ�.@-b�I�t�"������s�n���S�J��ՙ�<%ґ�e�x�Dy��T��V^�\��T�K/[q@��5��S���µ���;��{~�K��g�N�� �E&�����������:83X�,��i��!�L��=\�/�\vL�Liҗ#�w&x�f�$�S{ANL�'�_���.g��4�k�H;.��������`������l]�m0][�S6�uJ������8`X%�L�v�x�;���g������["�P��x/D�_��l�s�5C�͡ܪ o�v�[���};+���õ8�����7�΄��	z8yxpv�������H��U�H	zˊZ��D$����^C���0��7G =�z�y+6*�B��� �;F~[�IJ�W�b~���l����丙���g
C�2.f�G��k��b^_�1�2��EH�m{e��;n�Jx.����/�r�7]S9��MQ���G�DJ���S�}�����uT. a%|�����Y˪�ϼ�
$����@@f�[ތR���y�b�c2n�W����h�r`ĕ�X�>2O����OD$�!����������l8�a@FS��$�|d>�/�[<.�u�?`9ҧh>(�lṝw�Ҍ
�
`��F���~�͑Xڎ��]����bs��j�x��C���$cn&aVR��` ~�i�Z�R;N�r�t���ȣ�N�*�<�t����0b��7�Aݘ��Z���̨\�N ��BBTC�Qn���M�""0�J�!KTSam�����e��d�M�ua:��Is�0��#-���h�3{�&ݷ�"c4�s������Z�b���؎MmZ��`�&z��8Q{~K���=���|#��v�Gv�9+v�	�<�E�<
8m{�٦)ɘ=���Go	m��E%�Gͫk��.;k��W�!`�Ra�����v�
��yȥ8���.�̚�\��ߗ�@��>��Ł{ͯ�,;���6�dEX}8(b��)��_z�d�Z�,�&S^4z�C�4[���Ҿ �ƍY~��7��)�Ή�&��2��f��<����)���S�[��=����'4[�s���K�87��.�m��Uˬ��x-��C����x��3�[V��	Ɖ5~ذ^J;}��Œ�4S�h���Д���ܛ�U	NLw.����h���ݺ���P*�x$T�PB���p{
?�B�XR�<1�r��V��`NPo�ʓ۱w��EL陽�����������7w�P�M���F鸒r�J�hD�AK|5��ccڌ�A�P�/W�M�r$g_���c�W�,����$����z5� j�<1���GRPIM�WL�A`�Mv/*��$3�! t I��m*�R^�z�0�O��!״Q��7(�R�k��U�>Gd�\kU0���sb_3#1]J[v�U��.���n�|�͎ǋ�i��!w�	�~i.Fb���K#<'�Z�<�:��q}���a"�ˠ�\���o-2���O�1�@v:M�z|W�����D5	��u�!��#����JZ����|�M��]�`с@�YI紣ꉉ�vo5�.���H3�@>Bm�&�܏E�����&�	���6�bP�����g[�B���Q~2������w�5�]Z%�K��X�ۛ/�,���,��� ��r�RSv\��$*�h�Ҋ��Mx����G	ʹ�~2q2,4�P�{u�*)A���&-�De5$�{�b;��K�Rf�3k������^z@X0~�K���rث�S��*�B��z�'��|\[�=���>�(V��[��Uq)=s{8e�%�6�F�bA�,�#o-�����
|��|ܦ��~�2B�N!��W��7eFwb���Q�Ψ&O��Ag�7z����
��$L��ٻׅ�oI�wC؄R��5 |͈q���w�bB��Ǧ>D�]���ߓ4�$��9ay�����Z#l�^�S��mS��`��l5L�#0����g�˱�����"���u.�8Q��P R�?6�|3���
�P�=��Y�By����:bi�[O���2��t���O|ka�C}Ƞ�+1:�`����A��L��t��Z�38�zs�1v��Qm���K�T���Г���� @��Zv�km��R�A�Pa�dl 4��������D���d/�W�8�nP����N��֌�)s��C��/��M�ʝ,�7H4o����#��n5؋�7Q���FC����x�*>��eF�]GAiC�{5���H��Ϊ'�dy:�o6+Lگdƍ�0&*�Qyș�ny�:��T��-���H�A(����э�e��_\ �R�R�SbD�O'aj��������fC�ʊ�IP��=���T�3���%���j2-~�G�T)�N!��{#����aNgȇ"vl�>��n�~C��A��*���<QY�0��a��2R�زu�:���L�uZDU9�[Eĭ��V!�R�4N��̗nb�:�iyxD805+��hW-Pjp\��MU�	a%�rpCj7�[S����2����`3����BV�>���r��������{�2�n����F>UK��
%g��פj�1����
!�4
u��֍�K�t\_�{�z��[S�7��o8���Kyn�������H4 ʚV�W��ɷ{���tg5����J����A�1h�ц�����ww���~T����)ɠ$&p$�%[(��^bj���6�( x���6g�%X�Wt������b8F�bڏ砖CD*��Sf�ʣ5�[�v�zV���ީc�zHI�W������*	����{�l!�r{i�����������R b��@;�!<&�վ��� _m��5w�	ȿgu)�T�|��>��ݭ�o��MJ^���)�����T{�}��deK�yi���9��c_��Y�yD�PG�.3��Bu	u�6��~b������P��<�H/����=a���ź**|�'H��)��|�j	]X��������ՠG��& AbK�]���K �S��l�`xh�|�#t�HтH�se�փ��8xG���xQ�W���7�JDF���:�վ;���d͉���A� ��C���_����F�?����$������s�/�j�@n륺?5)���i��;�M_��"�!�ڰ�£/ŉ�����Չ�z R��W��۳U���\(%Unr-:͉t}Sϊ=�4"hTZ���(���b���~i!��tD@�ae�[k���U��"Å+��l;�j��Pʒ�Iʨ����8>����F7"�����i'�[q�Gʨ��pz�\Tj������P�Lg�cUR/�� �^�	E��8\02s���P: �7͵AM{��ԣ��u)���:�<�ӎ B�/ G<V0��<ؖ\&Y��'�s6\4� N���^Ԛֵ*�9����K�B딐��<RK�63ܝ��tڪ�LN&JI�~�@o c����Sfg�gqY��i��n[�CH���1���6�UN���� ���#\�$S~	��.�X�t]1pZ��0�ZҬ�,��]蛣��.f� ��-03c��$�,�E3C���=
��� �X�l���Y�^��J��4�to��&'��jJ��Q?x2̙q���S`�<N�=�M4ڒ6�._~������<�[)���FU ���;4}�� ��-�fn��s�
�!ϩp9�Z��:*�-�G��%O!w�eݜ�[P����5L��6��
^�A�����l
Th;����1u�`�Ͳ�)5	.��R��!:+~�s�Aa�����ＹY؊�E��7jH��)Ɲ-g�g}2v�sn1��B��`���8\��a��#ս�y��"͢{V���&+�d���Flf��j�Q����6��j!����bH?I�����L�z%G�훳�ۛ.@�H�p��.dG�v���%����X5��%vE�~�X������ڭiՒ2k�"<C?���H@ɝ'�@?��~`ir.@�i4��,
Er�������3����DI��1���M>�˫�a2��øa���\N��g��]`HbrS�r��kD�c�E1ƕ��"[�ɼ�քG�z���%1�|}f������D	He��txI_�p�����4�,�Y���_ُ����μ�%�f�gw9�f�R��
Z)oD�t������s�t^
h@����}F���`�Wf�.G�����Tu\���Xjy�v�7E dmM�-K$�]�_5���'�@�C��e�/3.�W���ң�	����_n�n��mhp� 	0�=hx�g�/�Z��E>��se�v��}:�R�Z�:ˍ;>���fgN�S�����9N����n�ٮm�� ��+��>Q�\T�{����!�K�\�����8�C]�Ep���u�H�tu\����+ڤh��{��Sfjl��[W'}1��캥�F�RGH���aEN�+A|l|Z��>�8�[�g�"��Z���l z/]�K�DV����
���mT\�kk�^��ӡ�k�T�y�^V�o�T�q���$�&Na��#)3\����`@l�oj,�:�֬c���v����Ɣ^����t[��,vf�J��'�H/Y�/�O!��<�z���jg4�lޱ�#�dZʦ��6?+r�|�WV� �����1oC��T�NpdO�}��P���1ިDMQ�0	�f9�>�ђ<fpЌ8�fn��!z�ʖ}�����zq��?~��;4���4=��Z�U^�i�lO�+��P���$��u0���G?5��p��I(|rLCƂ}R'���w���кt�?�.��Wiv��n�̑#IJH}�-��Ï�Q��i��a���=���E�K�e��h
�7HC��t�� qA_�ֽ��J$#����8��[�� .�H%T�
�qz�^H���p��T�$�T�i'���yI�^2\EIo���K�խ�ڧ����%�X\�,��i�o~�e�<8�ΥL�[��2~�I�B�@oO�1m�AlL�h�]q�?x�-orvQ7��_��u���P__9u#���I�p$v�����6x�á6�,>
`�R7V�D�q}9w�c���M4<,������
�Xb�*�b���/����kCZ~���t{��%�3zJ�&���?&�4\4��]U"��O�T�`����݅�����<Eq�G�Ž�P�=�䑮?����
����Gv`��N_����Z�3�e��-�	�U&ڌ�
����f�fӓ5�W�$��?�sH�,	����h�� pM�"9x���g��g�c0W�V֦���U"J:���=DŌ��D8l�{���=(�@t�=}ie��.��bq���O����
w#h�J��"3I��x� ^Ҥ���� �b�q����-����;Bs�:$��"(�Q�N՚�ู�x7muh�_��U&n�v�#&��˄����u��_��;�!�Zʓ&���u
ʛ��]�ZI����hX�%F$J�P�f�o�P&kb��I/��bc�9x�w~��+��B]�������}���nOh~Gan���~sF�D�{���/����x���Z��r�Hg����v��Y;����;G`GQW���!�<���� ��\���IئHCP)�nC4��d�J�:����y��`�U�Ȋ�����w*�Kkj�6�c�e�s��'O+s�0���Ǿ��9_�@�M�z ��@7�dP�N�(��r�(�N�nD�/�M{�w��jP�-��y��j�v2�K���mۜ 4v�SJU�Mǽl�����<��O���]Fv4��5,�N>T+)�kg�W%`��:�)��t`D^N�g��ocRl'xV���W�ż��uжU8@��f����R�&O�ˌYV�A�VQ�����bR�Ew�=t��=~琋���1���"��!�������p��L�J�@�hdլ�b�G穘k�Ш%J���DA��ɡ���}��?�b��<� L$��x�v�$�rpe�+���lcy�Jr�1K|�!���v����4?�F�{�U3�������[�N�otr��Ó�s�!�Ʊ�64V�.:����Ɂ[!8�X0�WRH�%g�d����Ʃ�Rv�m�����A����C/�M�6��T7��]#+Sb���a10;cqI��y�U%��C�ӕ<]�5�4Bh'�����j?���U�0 �h6���B��Llg�!y�G�l�"�4,/�{��Y%�X����/(�L�>	Q��yq�n�����6^�w�*�)s�PXKu΅���R>[{)��8e3ܕ�{��̳���Ǥ"��TC�J�pbt�أ�n&xE���F�R	\#�I�����혣X������,{����ܐ(xr��Ͷ��Y2@x�g4�y�S2Դ1�P�������8-��N/���j��pi��h3$�6� Y�/�,�:��H6���&/�0��ۍ89�&�H� W�I���l!����+�n��9��N}�=�yL㪨���:� >����0=#c�%rz��a@q�,�+�=]�T���&��O����l���1v��W�Mj� 	����R��د=$Άfw���&�N3]�J*��.�]����d���ݝm�$)3����$,�f:�*Pb���SC�1�5Ѕa��W����f��O�2˿�K�f3~|<x�+�xB��ǎ;Z>�,�}�͚�)��K�|;��֫��X����O��Q;��A��bB0�x1�L��&�XB=Uߊg�_dP��o��Y&`k��5.�����$TK�SVSsz"��(.�D�+de�3�4�{b�^h�j�D[	X;�t���]�4�P�o�h�&@k�6�h�V�B�kv�0S��֘�?�@9�~�S5=�-.qYŅs53�CX�L���YoSڂ�Ԡ�Q��̽dQ��Z9�f�z��у�)�O�rA�sh�u�nv��b�\O����nVpɴ'���k���W4Y�3\R]�.��QH���KN��sx?�o9�9@���93���"���>	8�幎��w �{�n��d�!|	�'Nv�W����׊�/�2nZH���8�3�JeJ�BN�,��h3��`|������a��)�q}%P��if1��L��@��8龓���ģA$�c٥�ٚ�J��n��*���͑�S�Ċ��?�F-t��5��Cϫ�j::�d��o���)���H%��׍`�&H�c<~��A䫀u����ش���bA�0?�3��h%�anl�H��2c�;����N��՟a�H�e�2�ak���d5�wl�pص:�[�B���fM��5�s��'Q�e���GD�Fs�����C#��������s�oު�= �1&�T���ص���G��t��ϟ�H�ek��m�:��@�:8�p�l��W���[$G�JcKaFW<FZ*�<�Q��')c
�/f�dK��gk`{7��X��Āa⢳�펬U>���MD���QE)Vs�p�R
@U_���F��@���fɬ���6�H\���}���;�4����*�9-ĵ3���.�0̽�����O��ł(H5|�EE.�����N�؅m������y�W6����XaN�i�S���[��.���C�,F��TYQy���T�M@�mf�
{HC|����U�����3���ٔ�<q��yK�+ԗh7��pj�7J�����xq�а��x�;6J�tdr<&���l����;�Q}\��	�e#ę���*��=���=�x��G����k�?�R���RW^Y��/��Ibo�Ӻ0]������0!��Lp�����+�-�<ו}��l�Q�	��� /H�6z6��A������Um ��4�c"�7\%n��xcOf�p�3x�$�M�;B���6���3{ќA�Zٝ7���=�<F4!���&v3gQ:D�-������G�TN/��っȿ�n��G����}5.ިD�Wy0$�:�O��=��3Q�k�܎�d����*��7�l�S�8�o�����ɲ�����r*?�w�f&��>��H��	�����d�&<`�Ap��F���ٺih�*/	�@0��w8Y�nK9gh�Ⱦ�陛\�hH�m���5��g��|M�i͎�Za����P+�]���+6w� ���
e�ǝ�Mw9��s>c�YϽ:�x�T.�
�y�*8F,�d�M@A��M������<�|�Q7�iR�+�ҹO���0�]f2551b���#^�9�K��v���?��{��I����=y낧bRܷ�d�
õ��&8��Qj�q�tb�"�� ;���7�M�}��ͭ�����۾�+�N�8��N5�^�Gl�M���P�L�~Z� ��&����v׹I�_��a���	�B,G��tFs2|�4|��l���[Û��ӊ.�9�;ܟ�t���z�7:�h[�*�t��Z���A���eO&W.��{դ�÷���kɊ���� Ȃ��OvEB���}ovs��iBS��?�_P��
�o;�xd{F�Lc�,BF�-CSu2�h�pc���Ĉ�1{X�U���|�#Sdoklp��t=	���6����a3"�C���{
��1;j<�������I�`P=���U_�<��`��������ғ��{�xTއ
���s�M�,��ʱ̼εP�2�Ѱ!�C5Ȩ�}gy""��^���:�Ϙ�3;Y�k<��QE�dwCOu��	�)�Y�C��iGO�Ӛ8�0�ۏ��R�J	L��9��Pd���t��"��������u#t�V����A��՗勒=���L	�k�����"_�L��¿�3�P�b���x!�`�+��#
�DD�6%�.>d��pa�`�8%"�M��Q� �
��Z�q~2�}A��q�&�K��q�h!ۣsN�!�x��P3���nC��M��ZCS��(Ѳ�'!��$����t�z��rf��"��Xax�ÌnY�$I0�۔����ª!}��/& ���;ɲ=I��HG�G�lO��/�D�h�gm�\v	ت!d�� ł-qzFZ	��A�i��T�HUCe��	~ϧ��~���vL���Ԑl�l����'6	8���~)�`�𫊯Q�RB��a�Rˉ'�c���ji��\�+��ò�μ�<���G�n�!¥p��}`��#,B�B��9I�1=��5�m�'�' 䩗 +H���0�̆��g-�R�K����������6?��z���J��J���Y<YfNk�?ہ���&�F�1�{����4a�ۇ1$��l^{X�G3����]�!��E��ƈ;Ȉ�ˊI���>=�oV'�M�T;#�}��l� ��sh]�Dd��M�!�HBf�5ꌥ�^R�koN� c<��aH�?��nL�dRH.:Z;q���P�������4�x���jߩ�(���j�fɤ�0�y��C
�u,,�������^D�#"���9`a��/H�g߃X['��s]�65݂��bU3��m�x�L :��JF(�@�_�Gr�y��:�3'A01ĥ��~�)�]۸��ʞ���"�B} �v�0rt��"��╧f�!)���KG�u힗Xv�v�mC*�u�C��+�a�d��*yY0d0I��7%8aac].�D�E�Y��{��5�Q�b��3��m���SPXv��!K`�V���e=[gDHS=c��n� t�n�$�{���O5Y�uoI���&?W��M7��?	�Vn�K<���{�v�Ud�߄t%,���<���$W<ϫŕh�~�N�R�F��!�p��������H���ve�1���zE`|*%H#��}ʌmr�5]���}���'y�J{�d������>��!� ���[:NI�@�t�2�ݢEq'yRH{p�e@�KQ�;9�N�|ٮi;+Eǣ���y����n���J�I�F���^*���%������>͛�(�EV�|��K�$t�G+啚*T�-��U��i���k����?(��Os=�)��M����c��2�G��ZC��7Lī��D�w9$c߲"�D���c�pW?�E�l��;;�Ȥ���W��b����W��Ok9Z�M����{��bg�U�g��q�J�J�j���]ϋ>$��n� `�.�ȼ?�{P2���Z��p+ׂ���s���D�R��6o��l}��w�Tm:.��=9'jr2����bi�b�X�?��.�{�)G��w�����֎��g�)6
�<������[���`6H��ߋ�2��%ǯp�|�6���׼�j'��6*��*���Lkpi W�C��O#��h��ՊU���S�2��k�C�
�)aޜ����@�zg�"\�qx����vI�W��şȖ]��G�E#������C��U��zv0�1�i?>���P}i;de�P���|g-t�����&V��)K&��|�|1��-&��Iߗ?��[	xL*W���`i��<UQ^#M�{��K�흒�Ӡ58&A�+Z�$�Q�	q[lW�
��I��j;��@�L�+d;��_����J����S��z�
ґ��A�o��YCYmU��������1�ߥ��[/�]κ�?w�M���e\v_*���.������b�2jv�Nb�C����2��&�Y�i�Fr4q�Ů��9�q�FE�A��_��O�����]�7��h��ƅ�ɻ��4zqʱV�$k,��$��rƺb�i�d�-v�h��r����VX�qǈ8��A}&-"y!�Vc�#�Y�si����HB����h���ix�~�-��{4dw�*�F����oo�`��MpR�z����	����>�78@x�Pk�<�m��5�� ra�ĥpi�I{��2�}2*��-DT��"��@H
c��eK�O@���_�0���[�8U/����5(�o��>��$�����2���FC�g�5Zχ2���rb�1M���&�G�e��;�q�_��L'i�N��}�̀��R�<K_���(�l�M������hB����li{˗0�O9��VMa��T>�����I9�!K���cj��n����]{�G~m%��"ĮYkҒ�E1�e��6�[+Ϋ�t��d�7?��c_A3�g:������c�n(p���{��K&)$�$��l�<������Yd���v�Oh^�.e
e�a��s%N��pI�mkU������
�Vz���,:�/Oe��ܤv@���_�'��`�s�y��=;�`��T$�F^������gW?�ݶ+���؀�h����e�s�/�M9�1��SA�q_����m����Q�0�@���yQ�*.�<�;�6�K��u$h�����ӼU�fS��2(wӂfH�G-ݢ�g̚�U�Q^EDt �@��"��t0u�T��K7k:
�U���$�v[���������F�r���	:�^��fPʰ�_�S�;럚�b�j���2f{��g���4t*r�����A�K7W,��c12�0� 
#��@�C�rA|
#~(w/�W�ݞS
�QdʨaI<��K5`�V�~��&5�U����7�k��Î,Z�5���T�OC����IpsͰ���`��_�}0s&��I��rQ�+}I���qd�QF�6��H�?����x���e��Π�U6*���.k�Y��l��	�!38p#�8I���ߢ5���J2mI˩Ӹ_�]�� ݽ��Dd�XR�g*%���K�O�:����,���"�����ZF�"<����^�^��~ʘ���S~�`�P�Ò����qfq�m��\��y�~��9�,�,�f��n��V����\,nUh�c��=]�՝$�k�tX�����0�Q/%�$�Vq�ZB�4Y� �B<��^�T eB(���RP��($���>m$B��HE&Ѕ��H eL�ȯ�N�[��]�թJz��4yT��5o��Dj�	�y�U͝���$�}E��6��w�<��֛e	���"�FZ=x�AIB���P��I�8 �h�Q,t
&��hʯ�}X9�>M����:N� ����Q��E��g$�R}�{WMd�3�z�#���{�aa��@�%7֕�����.�����S[�������񺯄��nUn �������Ѳ��E-�3���sܵ���1�Zg�a�\�����(�l	�-�]�H���`�B�&�:�|y���;�8�Vz������P"6>Oԃh��|�Wr|"ѝ���$�0~x�����uW��kk��D/ �p�R�m����t����\�-��%0&Z�"��o���T�����s���9�0|��*��"ITGK`s�P��4���HH�� 8F"�O���1�Rqh��?C�@Ї�"���8��}��y��v�|Ț���bʩ��b�O䗇}�'h�g�Ė:dz�}
.y��[��J����DwGB����ڰ-��/����TL}4��'� �}FD�r�{�[��,�w�:��w����u����<��a�� �Հ� D��Ss-HK��Q�X�a��<��o抔.�S��lt2��>"�?�8�ߋ!���iQwq	�V�k�A7p�ݲz�F�SA� %���;+?c��T�㺫�ѳz6!�f�1g��dE��P�5�� ����g8tJ�>���1���g�sX!a�]��루}���|{͖l��C?8_JZ_ق�Q�}���'�esI7Os���g�E��_�N�H!R�q�ScoL3q��a�Di��Ss�7��>�@������|�
���h�w�F�X�"q����4�v���)7��I��CV�bt��F����@n��.��6���4�w�U�E
}��\�uY�����|ޥ�V 9�H
��] U8c��4�@����³�<e{"]�{K�gp�5V���c�{�Ե�' {�ą�X&�j�E��-�9��R�Q~�gv��+@� ��'M}pQ�pͱwmz�s�6��8�yBU����wR�d]���&z�덋�������"�����!��2���jkV!�RqY��+h۴P�?��ߔ7�Ј�|U����P�y�*E ��a��f�OCuc03ps���.��e�.�K����D��*�r����G�:�e�>����P�5���Lc<L�@�d_s]�>���MH��v�;ŊR0+�S�2M�:E*�����m@���ءK�X$ަ�!=/2�����h�oA<�w��kUm�Բ�*3x�L�B�Ok�9���J�at-�Y�	ǫ[Lu6E�ĸ��!����b��_��L������H픢Gk��}͑�m��M\��[�6���;2\v�����FT��S���U.���%���;A?�	�ETI�+(fJ�«��g��o�#�sm� oZ9�$�:I�B�uh$k��@�j�&����µ<��_�фm�����\6�Y�#��-�6�ھ-r�{�zH�������2T���\J#٤sF���"ݶ�K��%p?�^k\���(�Wr+qMI�=�|����.pD��U�'�t�S����
�"t�ثD�^�#�)����l��5l��aY�-�e���4+�B��
uzΕ	���Ű�~vm�6M*8N���4+l����c�D��`khC��`���/����ۍ9`Cӄb_�Ľ�q�RS.C�j�����d`��%u�6�~I8�&Z�}^����"����C�;�E�@�J�Jm�����ݽia������nl�P�pv��_ �+�x�����2~�L>��������b��*�pX�����csc?�R5c=����������=Q�?���<�*t��A�)�t�*h��ڝc͌���.�U9��C&�d���ǆI
gܽU�&g�nC��'%P��z2�q&�t���*�]�?��3�c�a�R5=�dH-���h"�k��'뙖�]�[!b�9\zisK@|@�7c�����
�س?u7���!����bK`a�14�n$J91��9{�4����nY���ػ�Dg��\�$�׎ܲ��P�j���j���yK˴�㥏��Te.΢]��h^�v$vފ؞2ʁ���Z�a�ӊ:(2�YNH�6LT%~����נ��Cf��jB����*��Օ�P7|;JU���O��k��b���K������P��?u:�*�R�/<EoY�,�N�倧�nC�� hHS3��mr	a��m���sgC��"c��CXP<��S*-6+p
�j�hY7,��h�M�l���b߆�4ދ��'t�@zYu�D������@�)T2�S��f,�@�o�J3U�o��C[��PӖ@�0bK��;Y�����f�.DfyX���Xv#�V}�#�}��� ����	v�e�i������p��f��s�n摺Ҧ5�^Ύ��FRa��
�T`�;�|t�(X@�>���:������d���	�����'���R͕i��d��/��o�a�(��a����|��O>�70^����ǝ�!F�9�Ak�%)�P?-ۻ��m�f-nѹ�����|z�ѩHh�*@y��[�'���aη�9*�b�>�'�xiW�����z��aekPq�.v����/���h�G�Ɗ:gx&Z�E���]�u��M�6r8��5a� '�.����o$�h��#��E��ITv�3r
�d[�ە�����AM��9X����0kQB��Y�IUX8[5F)v~��i I�%u��[NfF�uc�<d=�V�w���$�F���h=ɿv�[x�MY�!�@��J�m���Nh9�g�5�������|f5)7�Y���K�Wش�w�o����ls���7�}\�*rTO�N�9v�YW�R�^�y�!>4Ò!Z��Ͱ�FK(�=Az�y�M�hbK�Ǣ�pz�c���^V�r�F\4�&��hҨ���ɵr�i��5q�Šb�T�Q�mA�{s^/*8��=YG%=���rl�B�?rה��zLc�aӇoB����]��q�cUgZ���3_
Q�~���d�N�<1X����o,p��e	4��b �9�����3n�$T&4M�����أ�7���	0��J������ r2���j�7����Xd�;�`]�?c�9p�)���U^Q|J�"(>EE�MyLP�?2V�?:L.��b󯔵�$�b�c��D�_�U�T=����F��(��4 ����'!�G8��ar����aL6h�xf�u�uoX߭�ou\X�\�"����.������\jso� �*M��-;O����7;�C�BX�dk`U:W��Tt�K�:v�޶����� �x�m��P���5w����pBS�;g8�5�B�L�9�J��xe�s�'�}s���l�c�f\�B-!�j)j�����???q�r��=70�^�5$E$8�n�D���5�p���EKQoT7$T��6
ir&���_*��Fy���=~�ZI|Ԭ'[��@��>��L�1�Xm�EQ�������s�?��y��� Tȥ-�|Q��U���3i�Ղ�f
=!ȼ����f����I����O�V�G쎷�yj�&�@�f=3��4����i�%A��#��y>��֑xQ@���n:X��㴨İ�U<{�{�q�@�U3_v��@�ʥ�o������{f�F�(�D��2Fc�Uf���F��R�_e����S/}7>Gt�H6�#�0`쏵��c{�|��s�5�Y���߈�aW�۱��	)�����`��2�dz�PJ���|!�g��M��PJ-�8����况H�J��3���O��@�"G�Z�z.���(u7$�5����®�Z:Ji;�2�w<��"g�lX� N���6��ʐ8K�r�N���Z��_�`?��;bbivT�
��?�Ly�^=8�V�6D�ڀ�,6"
��='��Q��
��a0���/���&	�!*�|��m�ul/Y�Pn<;�͘V�Cm��9Zl�M�A6�����W�"p�7���t� 4��\!3��Db���ˬ�H��ݧ{��(,�~�s�5>������B���`�|���5�k`3�/� ���p��Iu�?t����$S+kꩴ��8�Gr.����$�A/Ƿ8�`�5hj�9& X^}%��<gu*!�V��6���{8v��>q�#�h_�C���Y���sA��N�d�q�(�(d�A%�'�ڳ�[0���{��'����%�"��d{�1�s�ۮ5�P1m��\$}���-tՉ�T�d�_�o��	%��m1�F9K��Ǘ؎��?"���x����7Ruֱ7�ey8s��|U�!l1�� ��s��o��|H�D�J
l�3i��,[���f�=e�?��W ����E-�E��p;� �1E��������M�X"�WF���أ����0�^���):�B&��k�z�4�ce�U�j���)�i*��l#5�X	��ԛ��4�ǽꉐ#��C	�0��t��^��M&#�t�^���ah =���c}듥��\�m_�aY�l�\=�g��C`}Ty�����Aډ2�yzqƴ�/~hu��H%�B��>aL�<��h#�8���:��D �.��f�q��`�����TA�u��f��d���_��)Q�5��N���}�� nN���0I.�Hڃ�U&wa3��K�����Z��6�$
K�@ �:�/���Jք����E���芤�"<O'��8hb��W��<Qe�N�O��l?����$�B�?I��&*_���?T�o�G"�A�.TA����F�l�}g<��G�F���MO-{N�O�)����d��ԍ����)K���`�\��I��|C �������U��];etn�V3 �WG;�z[�~K��u�����}9���(�O��/ǰ�!u���:0	��q�W|��_l	]}[+tr�w\��'�1@����,�~��4͹�q��՟�IӬ��<:#5d9f�FS�.�!����(����ix��Xkw��T��z�>����k$)�d,X]>0� U�j�;�0XН5�E���PZ��P���S��}��JW �Q�LD��|Ƨ8�4/�#a�:������F��qg.cP(v�0 #|�8?dFhg]�?�t�ګ�,;���J�g�ǒ���ݨa,��/Ѝvxl�C%k%����\N��_kNuO���4D��ެx]�����$>AC�iR:k�����_��Pp��ȩ2�+�8�aN/���H��/�<W�U�*A��y�/~��k/�G��ͨ�&:�Ӄ+����:?�fSN���y�\��|��uC���Al��H���p�,v�5�Yr���\A$���(=��f�c=ᆾ�'��<��H�Kt�l�jUJ6���T�BT�3&q̓,ڣ�y��-&���
 a��.p.Cb+�����x��r���Z9$�`أ=F�����6ղ�W�&��N
I�kT�����Ģ$�l� Z�)X5����k_��!%e#��^V��G��S����g��J;�u[�0�"G�Y���g�jp;�,u�����'u�;3o6Dѵ����g��F���́�c'~(H-V~�:��bf�:x�(� |i#��T%h-��@[��q/�%�����BMvK���6j��nnW�ǫ��Lf��l2��z4|��X)��_�W�/�g� r����{+����=��Fr�^�kT5�����`�l��8Bx{�)
?��@��?/�a���2κ�ec�0ʓ�E�O�j����1�{��y�R�nR��i?�D�[� ��C�$�DP|�0v_�ƈ��:G&�1�%��< e=���p�)Agw|��ާ�K����f_QK������ �=!���&Q[Ϧ�p��TUa�Ԗv}FC����ʓ��9���]�+p�a�c�T5Vt��5��j�X�1:�aШdd�?Hg�$6������f�~��.�i�����=��Uejo���=��	��{���a2���Mnw�L]��j�����p��DŃ�D���j~t�t=�+��4 �ZtJ'[��$�FRC/??yA`�Bq������P����s�q'�{ñ�*&����c��5��N�}:h�T�n��qKl�s�(Y��KS����+�@U���ψ���B2�JC30&�-<��i��L���l���,��F^0��T@�> � �	�ҫ���-�/T��������S�]�U+L��Mg��pIh��m�Y"����K�?������\nCs�N�%�[��S��Ӭ�7~q2��WYŮ��r���U��߯��ݚ��JLN%����0J�g��hS4Ʌ��3|��.�4E�K�mߪ����JPP��.�KjO�(�
}k��B{�>�P����C��_e�a���H�	/�h�R�)n�0����Y�7�����%rڢ�/i�Y�<n1�I��gһ!{�U�0���S���^�;<�C�1쇫M��^�N��Z~K{k��j׶D�����d4��f�lt�j;����$hT�6��}l�C��ֿ���(�:M��1�/�N�!Q�L�����u S�xH]����ˍ'�C\%�l����Ȝ���x�P��z��!�a�B��T���O.i�@,ǅ�3��Q�0gId�Lƨ����JZ���u~|�v��wJ�U�+�����u.�cI	u��Mr$`�#�Hy;gUc�*��a.����2��oMM��N1����0�Y	��])�����G��߰�Ox�&!�$[��1������\�oQs��qӛu�x�������" ?@�f{�������!�O\�.�G_�Y�zb�1�::Z�#=�T�(]J�DP,��������.D�i���&�&��
�xxK;jf)zPu~���3��M��8���+'b$�Ċe�6谪lՖ���y��%����9��L��rT.��l�Ή�+6S��=#�"�ɼ�ߍ��AQψb�J;\?_ܷ�.�Ś}�	��RYA&v��~�"��)�.M�L>�k.7DS��04n�����ܝ��C�d�#Jc\_4 �5�*�{ص	��x_̱"1yT8Ǩ	����0�,^H�tH��CaE��+�|M��2P��2�k�b�RQ�X�y�%����Ga���83�j�#>�rz˿�?k���\��ޕZK�L�	h�%�u�W���_��dz����p�)����:`�s.�"Z!��93��[���%6����6�v�#>1�"��O�yx?��(�8H�Bnm�Y?g#�c9�*{B�U��n�,�O<��eڌ�;MW��D�f4�Gt/e_�k߰�cL�S�eC�eI����3��(\;�w,̔�n����/t�{Y��ħ�^�S��o�+���$��|�X�
k�~K kR���_��	�<a�?��]�SY:w%-�7w�?��9�M?3��d$���I���Ã��c�H��h�M��gG��k$�2t��:�5~�F�AjX(���2ɶ.��C�㦑i�Fu~^q�SA&�����(�J�5`�rV�!0���P|dw:��  �x���/#y���5"Z���m�ͣqu��c|Ѯ�۞���⦾��N��L��&o8��]�TǸ&@�$Ӈ�M$2�֎�Y���w� �	t
��| ��*���W����綉m�����w|��� �W���Rެ)����@bo�6�Ǐ��o9mV!]�z�@��ᢃ�c0.�$�K�͟����F �L�K8�®+�)]S�����h��*|ѐ�>����\�"Z!f*mԐ��x�/�zxGE=�//c�&b�~���`�� ǫ��/Y�>_r���H���+7�����+1n���y�0\�@#DIԮ��U�v���!���ă���z.}ibşS����:S���wHxZ�:B�藋�hQ�������x�L��ԗ�ϙ˹�{C� �j�����-,�h��0.�e2�=W��y&C�a�k
g(�;�モ2�wv�uP%cud[Z��pӅ3<A�	-\5���碩�*�����1a�S�חL�/u��g�Y�C9�FI8�,cF���~7i��n��?�(��]�9~��B��1��X��G��S@��mY��ouH=	�&�=��1�6��K���j�P�}��M�h��ųC:�P����ֵV��I���W��LĆ�"<���rQs;�������b�X.a�����D����Ç�=ĶB�n%�\%/�8&r	�W6�{��4�Tڕ{wBɹd[jV���7,�GP�_<*�I�h���r}�9���fLOZAZۥK���w.������^�l7S�3�*�`֖�=U ��6�	��bZZ�D���aFTyԺ�,ǰajs��p��_�?y���<?��|�v�'\J?��9��g��k�7��wӊ�`��(+ձ�����ʰ��y���T�_:�IH��p$�w� }]��=�%����H�-���Ι���P�<:���=ae��xQ�%RY�-)�����M,�V��i+���@@W���E�ȭTX 7�5rL��[`���B�jx�cХ�ʮ��͖`�jP������lw<�����sL�)��5�
-�2��i��3�V�qgP�-%�����ES�!L�ƿ;h���Y}q���0
;��M��@2�^�r�U��qz�"akN+�p��;��� I�a)�������+����x�k?�Q3d�͊��IaƲ�$�3�K����$?�ל?P�9����ϡ�v��B���^̉��'����P޼F�#�г����ۨ�� ְ�H ������[k�≅T�}o���T}#Y��L01�v4��Z�`xM����.��m�'>P-/F����&�����nN�sNq�~�;��ϣh�x�a��n5�x2�~�%�=� ��$�Ԅ��Xh�Pd�*�5I�IcPs0���g�(�l���,P���2,Ң�R��r�-���[�}��l<\�@9���T��:�K��k��y���Bp��.5g�Tec�2B��v�}��x���{�pk��,�����	`�w)����08�T�ʈ�0�E/5�\��a�`�H���I��*?O0��d!�<|q�㶽�$l�f�b��.I�0�kƍ���M��4�DYOj�2�b��ܹi�h�jJ�k�#�߇�E	�%n�*'�<c�t��E)�j&b^UK�
f,�9�g{�g��u������ ����Ռ�^��d��Q�9�#`n��S(��R�T��~SO.Vy���.\��Ѯ����z�b��T6'�/��E��٧�|W��p���c�
��߭�4�c/@R��_$�B}�&���t ��2vӏ3a������`�xI�r�.�<s����G7>�B_�J�/���O�Y�31�]���%���:)�Zx���ݫ�m����5/ww��Q.
t�Z��u�Lʶ�4�LKw�9�F ��٦�F�Ҕ,(ˏ���y�ub��*�mO>	yn6��o��4�3���C�(D7(Mͧ�p���`m���S9.e�F�S>����^0a7���o��feW���3��v���yI�hcJ��~�D�����n���r�q;8D�Uَ�:
�ݤ��u*Y�<&[%�I'���a�ըף}�W�S�	�)���}ѵ�vxZ� ��,�^bV�����&����������������ƽ2˝��%4[�4�x����#]u}
������0�`�E<+��L���hk��U&�uz�2'����M����p��K£q<%!�3�J��g\��o�ZD��dl�ܲI�;��q���D�;���.d�������Q��T�Y����w{���E���u��!i��T����J�"��<b`�H�5��Yeך�!g;$�ʭ�A,#�'��,�*�k(igi�&�VU�o��r�uW/P?�+�Q�M;u�Ǿ�7;��wm1�%g�
�����ͻ�Lđ�e���u���P�I�L�[��Y'l�d٪�*�b���g�s^x���3�Y6�?	��rA�̠�Q�y�ꙣHa+���B�/[��?�;�L<$�>s��D�5�U������\�an}�?��sf���pM��A?���9�z8�@�N��]���HT��ê�d��%r��N��yz���Rg=p)����w���{I��Q�����#Ԝ����/@��+��(:�J�evtش�U�$�C��2v������x����ep*�W�J}ꪜ��٭e2A"�"���e�?8�W7�. /)��ju�8���ۨ�["�ǠZ�]'t�Wxˇ��X�S��9sw�/��k��hQ�sb>�5���nm�#b�e��h-y9�|��+�	XpD��)|���2��siKZ��i\5��b� �&4��'3��r��T��`L�90fU��2�\[�稈\���*�0S�����u(G�U��ҕ�x��{�E}��wlޚX�BX��Gr1^L�Fr��o���s{5'ͅ���x����f��䰊p�M�u�<�;	��͍ p>�q�Y���<*k���|}.s�7�O0\(iB�M>{_���'Y���k��F�)��V�6�����tx��d��Fݞ]CZ�ĺ]�AKX@���'S�)���t���:c��.�*(u�U����Rk�B���s
8�!�� �eqx�Ce#�������q:�岀�6U5u_�5+e�ٝ��=�9�2�ks;.C�boP	���0 �_	v@ܳ3c��g
k,xҸ dF��;r����,�:#��3 E����(�� �L��h�8������1c��>6��ٟM�r��j��5�'���B�1"�Ö4��0����iE	��^N�\y���p٨	À24a�*lO��e������]��L�exm@�{���v�m`�sXM�$c��~� ���նv��٣�8�G�'6Ў������U��0'߆�m����i���|r�'l��{�?g��´���!�f�-����nL≩ˆy�J}A���p�G���O;����H���!o?O�NYǾ[$[��d�l�6Ƞ4� ;?�/��`_DRi� ��"�I)�o�mY=���<���^e�ĉ�t4Q*��a3g�@�N��[AE�-����C)h�ȼa�9	��z�c�i��ӛ}T��VYu�b�X=�x֞˵7$�~i��S�Nء7����]�����˴c}i�(I�fj��	�x	D�\�VJ�o��,��\]�6H�;wI0���̺����x�XjW��������K����V�6� ��5�yb�2v�Ye=H�Dt:�l`�ؖm�\��Г(��OM�g��u�>�s}���T��%>��Vi����w%M��{}��,5w��

�=��+�+qHʷ����D$�����.P=1��]�4����-�kUX�0��I��ɋk�@�U;��0�����^���#�x`��N��?yRz��%�/|I'�mҷUo���w��O�,S ������}}�B2��%,�	9]�*�D�<��\-<x�%A	�LW�	47�$;Q6ÍE�9P�~���j�7��ֺ��b�ipKp޼���<Y��i�h��6,��hs��z��b�5N0�t��R�Y
��o�a,�-O�p�׼�JZ��#��k�&��W��AY?�Q��ѵ`��:'�\��|���-3	� ؆-͒)��<�˰�tr�Y�-��K����2�1q�O�%�Q�ş�BJ�x��̱z�@�O[(��qW�g��9�dza�}�GՉSX)./bk)a�AZ`7��P{�:����HK+�q[䛄�7�����{�� �ѯW��'xM�i���WB�,#b^F�@��+�o�<̲���Z�!�	ux�PZ���*��}�[Dٽ"/�{���Dy��$�Դ5F!7[9��;��*g��n��?����pO�sQ��4����Cb!�ƞ�O�#�2�G�� q�\�B�27�B-�ҕ[�O����tlF�����A�a�b/V�0���#���疝��^=`N0p��$7�&g�P^��_���mR�\���UC�3FL;�.Ɗ7���v&�a��P� X���U�����z�+��;�U5	��y�(�-�:�0�~�F�,N)���%�M w~pDW���D��xD$p�z��������K���2!�hDú%����B���Ib� �'�<S�-s��8������^ݳ [���qS�zݙ�� �C�a��@G��?�>ޏ�գ���;iVդy��;$&m�z�b�����ǵ�ƿ<A��x��6���R�1z\.N�ߎ�H���=����cRlo����v�f;�cZ�+��
W��FN�JɊE���s�'�Io�+�>����T���M��>p]�����`�it��>�0��zn���&vZ�����CK����ٷ5����!2A?0E<�J�_Wm4g|��L0*��}�ᷙ��h/ ������w=����`enAܘ	���Hsìp@>ҲA����J��K��I� B��[���W#^�3.Ӓ|�|\�*��)ՙ��.&@�����
���ϯN��A���]9)������(ݟ���-�vM
�ݠ�q�
�]IY��$��Qx9�׻��v�=���Ԭ�^œ��R0٣�X��}ص=���[jYӳ�|�4H�^[����t�p;�͜}�@[�D��|qv1x7Gm+n�t��� ��w�W��N(�O��ϓګG�����kZ�gT����a����K�<�ZF�Rx8q*T#� �jr$@�P[1��?�����A�!�����X��&'�5�'���+j'�Ģ���ӛe���76��9�e��%G����zi����~�L2o��K�{>.��vWE�p�MY��
Z-�}��A��E%FA�`P��&�V>�b������IG�p3,����&�7�С2_`�F�
|�����bX��P��XH���#�mؐ)��h�h�9�c"����h�d���n��[��IVyK���NX
>-B�A�B^_��(��[���ex�Ӭ�z/�J M9��~7���g99�f�yV%�N����:�Q�\OG�2	2�[�w5g�V!46�.
T�5���x3 ��aG˼�p��p����^����� �ҰA�AwRNj ��_�΅1�+6L�W������a�{[�*
�$�e��j�zY-��DX<]2�"8a��nJMnh�7E��מ�saTS+ ?�;�ҪN��V���?�l
� o^�[�	�Ɔ��( @�r����AW�i�Y4��}Ov���ϣfqa��<Z�'��L%��aG)�<�VW��K('�bJaI�z2��J(G~��
h�����ȁ��B�������M_��I���p����h��̀QSx�|�3�v�uG�%��\���#���Aش�b�K�z���G;��Еט�*��Jk/Y�#k���iX朧ZC��?� �bA��R�� �VE�O��ݍט���	$��B{@S��N�#oq/��qdf�W�5ta̸�� ?���A�KrݢH�d��-9�j
��K�?;���&yu>J�;�����몂����Y�C]zcV���7z��.�/ZV�t��p#anI�9<b!�ߕ���$Tv�V�Zظ����1zt���`O�.�4���U�h�	��[�N����K�{i�G���'��K��s��Gs$=�� ;yM��p��}�˞���!�i֟�pϵ鷈���{5�j�Mv��yh����G��)^�[ �׋&�[���MP�=�Ǹ~o����n$��F>�f�G-E�dL������2Z	c���*�L_���+@g�����䀏����n�@m��7�T�z>b�<z��O�B>�WW%�b����_*���@�*�g������K'zOJڎ�́�V(I���2(Ș�w��
D������༘a�s�h���w0���&��}FDS��PƄ�dO���� �n��B)�	F����b,����qB��+����*\��$�>���PY5?�i�|G�S�եg�Y7��y[���21���d�`����
��Ck9�sM�p��O۷]
.�� ��db{[0�P��SH�~H%R�6��=��g�X�"Wm�؛�h�~%��&�U鱻3>"
[�����}|�*��i�����ů.є��ߏ���g'[:2����>�[�P(�6YMou�pD�lʘ�~��쳐9�����I{ٺVy����0)=�s��c�,�0˨K��@�.碭m1k3����J7B%�WT8��m�<��T�u�h�eb���^����f,O}���c��6�ޗ0�U4��%*8s�4~���b�h�]�O�ECС���O�G��PxEA��t��	^���:�����s)K���5A�������Y�x6��1	�w�gJ%*�j�3�"Y�����"~H����	�]��&�
��M>���6{�ݝ���u��j�8ULw���N�tM�6�!b׉��#c>_0Vch�[`�z�8��ݠ�}�܇$׶�p٠���+�y�M�{��#���Ϲ�?b�MϽ蘟�Ogl..�10�!)I��U[�v)b���_�9��j=+6[)hh��.!��xo;�~ϞXZ`�xU=�y�Q���mK<u��E���]�b�S�e��$?�f���vt�
nXa�I���"Q��ov0�M-���g��6$�l�8�L	�~�n�x�4�Y�6��g��}dJΪ��7�2ݪ�|���Xv:KZ7
}n3r��Z�2a��&�T�z�Y�m�"c~���-��O[�����s��~���G#r�V=���9��8]�J?�?hk��Dh+0 ��M�� �'��j��iA�D1Dm8�Ol��z4؈[�Z��γ	p�j�Y�����
?J�@>u@C��5-O�L-�f��i��Ŝ6*8�I��GW`wwK/�����(���O}�A ���.�1�Y	�g" �GOl���wvS���=}�}�=iص�y�:����V�����"�/��ͼ�=���+�~���rzi�S�=����D�I�=Z0h�nҳ�-�˥%i��v��|cZ��Ǹ���t5 \���$���i�#IPۓKj����U���A�2�����_���#C�L�_����A���������`���^�Rɞ���^;R��u=������v>ro,d��� � ��V�U�m�ӎbh[��mY�>%�Q3�3�k�����<*�?0&��H��#&�^�R��iO^z�9_k4�e+��X,�p.��<���#��b4����$:^U�NC����Ǵ�+#����Y'��‹R-��A�x��%5�/Px�rF�/و�|��gD�#���Y�G �X�`�𭕓� տ?7VsNUx��)�%�d��ܐ#��L;:��\���k0k����#w����RIYܮHf9zi&��W��ꍼ�j}禶2ƅ�ȍx��Ol��:'"&Ff2�I��M`����w���7����{W
q��KJ�ГꞘ��w�4�av�Ց�W�md�N���h�����DA$`��v+��p���ȑ+q��>K���A�.$�D����=Y'�Ry��_��iT<��������[���~�1���*ko��6��FDi@~Xմ�X6�SnhT�d.�KJi����ο��
��m���u�Q/{�����D),o����x�x.8׀����`���P�x��a����o����uK���h��w̏,�=����.��V��"�Z�̔�g�ghZfG��Ic��^u���� �;ʓi���	=�|�P�0�\��F�P	��"$�C{�/y[%��/{�1L�j�G��O^<�P���ML^ʆ�z�]������;�����h=vt�z&���	���J:Q˱���f���j����
WWt�	���nl�	G*�N=Uzp6�KS��3A����B���`�g2��K�0�T�X<:��ɕ�s��ł����{�zٓ��y�]�d�m�	��&ʏXUX����Њ�a
b��$��αDF���&j�
�0*�3mp�'3J�* KV�_��r�ְ� ;J�S;��>L{��xq7t�K��9g����u�X8�Ml ����cٶ��L6��hwT�&��Ys@�ڝF�"��@Z4��3ߐ�"i��ܙ@������wT}uA x�>YB�@!�y�FL��(|x�ҳ�w�&ـ�q?c�S*�BĻ�Hn7�:a��� ����A8��m�ɜ"�|/Ia6ܟ����}�M=VA0�R�C�/B�o)t3:�uO;�TC_m�냣��	i�۴H3�q x��V��d�L֔�ٶ��~q���>g{;-qݩX�أ�|!DЭE�={���ބq�L���mkG@j�q�����y���)S�SJJ3�b�=�P�P��W��E�~����:���k�p��"���&��LZ�;�����v��f����x�@z)�"�u>���M)D	r���Jw{d^p�G�y�5avI�(䟭���x��3��>���2�:�7�q�~zw���\�O���E]?dB���V���07�����
�p������ pb�@�
RO��Y����B���� Ԍ�oH�jCÔ�N�	m�D^�8�w�2�Pw��n�����v�}g�D�!�?*�:;a[�jI�|4�	�l�G�hm�KO����M����k�@�yG�,����4&zF9��'=W�D�W�J�x�;�K���}s#�qg��F�NY��>Y$.Fr�g�IGc�T���]�VwB�B�1���ö!�}D޷�f�Ղ�����S
�]缰!��1�0
�-�����01�����ĝ�q��3p���y'��bz�T9x_��Qp�������!Y�NK�5��j��賌N�Dw䏥>�����*Q���ݝ��X֕�9�$�*�5F���%t���-���b~����![G�nOl_՘�"i��t��č����U����u^���1/N'��7�u!���6�{�j.þ]g�A�N�2�Y�ߊ�+/��h!Hb�5�
W�w��#�9��I95��D�ܒZ�o	�+"�:��S8����+����e�Jf��PH��X�S�,�q��Wp��Ȫ�M��fk�)�p:�����@�#��.Q)�R��]�e�C�1mb/ü��]�p���z��A��*�3�8�eC�1�V�d��\�m�Ծ�\�_s��W��.t�m�W�g'�U��~��R3?�(��3�s;�"AFV0�#�f��g��p�Q� J3A�-3KM%֫} "�6�¾N<�!Waε?��`fMح�%�vѤ4{s�s_��P����b/\�R�v�@��e˽��WN�C֋���0נ��ϵ~Y�����:�aI�`���h�or�%���3�]-b��G=�mr���+�Ĕz�������1@T��2fry���e4���Ԭ�2&٩��7r�cR��3o��b��(�_����>��ؾ��n���P�\Z����,<v�T.v{��:��ɺg���k�$H���C�����R:��}oP�b�\ˊ�珝zH(�cK�/Բ=��o��:O��X$ԑ��X-[��R�:�V������U�иez���az7�=#��/��N�q�R�����S@���e]�u5Ē�����c��	w�I�D]i����ѹ�R!~,�,\�e� ��B������2�xZ!xDhՑ�ϭ�s�+��� �w���G�~�Cb�>գ*�	溯�Ӿ
P�'OV������Cҹ&��0�`�&�xo��;�
'���M�}���lȘg�Ё�g��] ������C�c�
tN7gV��"��$^Y+�Oc�������M�a��L"N["p�x6��ع\�;<Lsz������Il��4��`�d����/̸d�����V:�u��~΃NVC�P��`���%��J�KH �CS�I�u{T�$�ΪF�)�5�(w�xs��alR�x�MyX_OTL�s�d�m�.G�+F�m�ч��Ί���v!pn"�]�P{f��1t����zG��G>@I�15��Y�����YsߎC��C=��Y��e���8f���J-A�+�>?ƌۇ>S�Ɲ2º	���y��0�n���}e�n�yB�@�Y���S�2`���oN������x?D·3�k�6��i��~�yuy?��8�(����c�F�EW�o���-&�qp7���ڢ���S2��%��=��˘�F�6HP���#u� $Lu@�I�Z���y:%�����#��ٱ#j
�ډo�ꂤ�D��l����_�1��jvF���y��w�����Y��i��Vˁ��_dT�*�,��/��U�%xQ7�>!>�>𤔳?�fmy�<��HWB��a ��w��O�b)#�'+��o����;}<4�к��Ł��@î���ѽz�8�T\WL�ˬ{���q����	ذN�/�6λR: �a\ ��|�#Qs�y�0����ȵU/�%6x�떮�R��?�+�t�㿭��d����܅�����ok !j9��a6+m�@2	��'`�-8|G�<���ʧ��qn/₥�=6�Ƭ�*TU����
&��S��`o��U�線���������q�ׇ�D^��f�*�A9���0���/��|#����=_��hC�Rߌ��G���p�d\�H��_8.�$��\y`1Xi�~�MV��a+��k��\�@�̕��DB����lb���0��j-y��ޔ�����N��Ч�OI"�9�?�Y������������C}�9,-��J��(�o��W��Ћ�r���q��!�C���e�+�0n-��=��R�[�*�fe�v��~-���R��_�2�v��3����x�Xd'�v>�� �n:���A�3��F^���BN�	"��9u�o���J�L�܂��Y���j+�
i�	������U/Ts�R�{�W�|~���\#��#��.|��pBRM��O��F�	��wI��]��@ԟh�E��ńc�m��p�#�c+��̮�s�x������I��cEӨ�""s� ��[�#�)���w9��7�#(j�5�9��)N�8��8�r〉�|�1ӭ�oǪ���9��/-�p5}���jĢe��y�I�wz�/�R:����8���2�2F��|��1|K�(�w7�JgsEG�K�p�������u���NH��mo�L��f*�x ��YR	���ix�m�X�_��j
�i�dqSWs�J3��dщ�0a��MW�	����,q�0���W>��H5�)�ݫ�P�:�/�2\���.��C?���G�o�p`_�x��Y�0������d'�V���C%�N��BoBH���9��Z2�*��	Co�f(�s�{u��d�;v�cN�A��0̻���l���ލ�X�\��F��&R���
���W1",�W��f;�ߕR���РϧeSW�g�x�Lӎ���{|?�	4��^5�g�mnbV���m$ʴR��'�^ܷG�M��s1����k�&�+�-wr�9A�J�������D`z��07AX���;�B��d�{�/S��|B��ISsh	[��ڛ<�Ѽ����掟I�'UP4!5O�V ���Z<	��r�͢w�0X��X�0�4�|gcu@����A�=�Ꟈ��)_W��r����͠-O�������q8QlݫS����*1�ܕe!{UHG iF�P������3m��������`�]Y޵_�s��	!�FQ&���Ԣv���C'���B'�����u`X��h��媺��V��G�ˠ`0�ɱ��c�"��6<�hx������y֙# {q�]�w���_��PG-�B�Y�s=U����E���
t+��W��q9�L��j�٨\��@�����3���(��yu$Kv�t�'�.�t�J�<ٶ�8�C�j���N�N����-�T�BgEh���w<����ɲ��d�;Y��y��Ş3���'��%�A���ބ)S��T��R�YU�Gc��n(@�r-���m�����wZ�U.t$l�*imJ*a�~Аv�0�����i��Y�� �*�U�m
?���Fq
4�2����.��P����	'r��V y���#k\�[ �~����{���z��,~�Ud��������,= fWŅK�n{X�lB�����y�IW�}�Ds�>_'Fd�tlC��c�V���e$i��?��^bt��9گ���߲Y0[���T;ka�0���]Dk�v���ؽB����q�C����JX�ZT�T�8 �5��u�5���k�S�P��O۫f-\Y�N�L�F�=��"��7���Z�Uk�5�@���*��z���Bmܺ�!1��r�\z�l�>*�(��H�->�]��z9f@L�g��y��ҷ���j{�o�MD5 ~�0�
����ۀ�����Vj�#ᙼCtY��T_׊��)vI��`�$�97w`��z��	���Ф����j0%�	����M0����v�q�4�g�'�Tx2.��^�ؠ��e݉l������ԪdVx����`��Њ�/�ȑt����<Gѱ�,6��=���pv$�d���X�V�O��
>̑?6��Qf{������G5�8j�d ��t��������.�!H�k3����D�wo�vzI]�U��\vU��c4����F� ��?����}M)�Q���O�)'mp�#���1�����캯	�c'���8V��D�Z}���[-�2�λ:#�,�4���r�fC�jDӋAK��ݳg(p@!e���!�{�5��wo��g:�����¯�xT��m�l��T
u�C�$��)m"������.1�����}�Y��:��e/��}M�WG�I�2B)풚�����[�����{��֊�ܸG+ܻq����/���Y�p��q���6����\dg�u�5H7n�5��U;�F~0R9Cߩ)�����P\�&$�}j�fОk��*	ɵ/�T��xEށ��}7uzґ0%g��4n��IP�y����0�6`�ԵmL���)\j;`�|��:�f�ҡ��:'�qW2D	�9�=�S�TmՁa����ܓ|�D����>�>A�6�^A>ZC�4��������<M�'�z���i C�'���2�ܧ��?�Fg�XZ���_lPﾫ�ʨd�H�VK�b�@`�-9UD�Ӵ���{-�)�A��P4�,�>��բ���K	� ��T���?rǜ�{"N���А�lx�X��$ɎXj	J��wF��GH[�r����?%��t���nd�����{A��M|�v���J�&��B+���vf�P� ��"v��@m��䗱�%Eda=D{��`�W�kD��6�$�̵��3#� ���ą;�Qy��0�_�,:�sowV���wg�	������qk`!hf2���6�&�R|�5E��즨5�}�;�ݡ>�Q�/"yԙ�>���U'B�ܱ6
��.��xA钎_��}4��y�#�w�,�k9B�^�ߨ
^EY�MJh�Z���D��	�/��&����y�0�S�h�`����eo�hkҖ&{���4�����}KPx��4#�z"��px��p�&p�
����`�?�s�DLdb�ɚ��p��b;2�պ�O�D!�z��}@"�<2�zMO"�H9p�gX�d@�?���,�=2�}� �s�* O��Q��`�D��"��zayro0N�a%��Ԑyf�Dh`�I��TY�f8�9HK��l��
���A��oL0����8�^�K��!���E�P{�i���
� �kz6�tӺ�����Huw���o�Ō�����J��CjR��s"c��-w���p�4-�͉bEFVxe��|(d��)�>Z����8�cC���,���2N���T��U�[7r����j-hO7��F����MM���RY�� c�ʣ�3T"�<7`���æ[��+/�� �����ߛ��W�6����h��6�iH�繀��'��%Lx�`��546���U�Tǁ�e2s��'8���
���|*��o�3R�0uM�U|zǛ�5�JOOzG5;�z��y�ar��8�캓�[2n��sӚ�k�E����s�<�c,)!q�;�ت�*}[j�����?��x�VkIB�6�B�M^�[�&���Z��"	���t�JZ��d#�|���&��gk�9@)��C&>�����ɻQ�ɧ��1��D�Tɝ��id�#�)��-D9(��L�r�i�?q�R���H���%5�9��!�y�[Ӓ4����4p��.�.��^�KZOp�:�Q|@�m���k[׸k���T!F�:zo�m�v���������ZC-X���f��f��g#t�$v�"!:L�A~TI��(I�uf̴���g ʦr�״w��l_~������!'Ц'ɩt�j�+l��-W��:?C�O�U���+��h��q�Q��6�=bA4_���G�ρ�ʣ��6�_�	#���aBq���#`R]W�ᵸ�����Mq�2�ў�?@9J��D�a%��8��!b���	d��gHJ�>��/�d�v|���}U  ������E�v�a�e�����7��$�Z%^��s����.��˺�b2g��:���m�,��DRh3i�q8��W�_q�Ez�S�l��ɐ���6��ȅJ"uyV��SȽ{���	�y�{�M|�l*��6%-�th@L}��R*4�[r}\���u3Y㵃�����a������QC�$�k�_А�V������#k��w)�)��G��p�;v��_@��.DF�R��M�_���f�⒨�g�u��'Rut^zm��dDbH���Ng�_�bPE�&e�]-I�Ӊ��M<B�̉Lp6����%!�YSg�3�\�%���z�7Fؒ_�ҁ�c��/j����Y�-+q2���=�S�Ai7=X�.�6���x��s\7l�m��
�Y�&+�UX� ��=SB����,!�o*��|z�8�K�%ݑ	���B
d4@��	5̼�*�g�j@$�������n�c��5)�Ճ�(ơgś�T� @����+<9r��n)�?p�ʰ�ލ;���HN�L�OO�[<��={|�`FEΫ@��m9N���is3���4[{g+������dr�r�/�WI�!�$�aJ(�6��8��n��(�$?�/҈��mӌ��J��Ee4u`�w�D9�s �=����^	�3A�8�+�����߃�2�ɞ���U1��w�X�bq@��:�OWW;�-n�K�AmJ����*;8H.m��O�h�IC��m��
0��%�����Y��b��!p1a��B�RJ����ey��|n�Eoy}W5�t-�m=.�Ea�꺷Q�A���+'oT�<S z#�-�ާ�q�1)���S���L%Q���%�!�>7���[aR���8-�F�U�	�S�߉FP4��R��*(��;�Yi�i�ǂ������6J�lb�����W�`z�UqN�{#w_	�,�� s���k;���}���!qU؋�&�U<v����f����A��.|�v����z@(��7�ǌ��k�`E�R��vKa;��s���+(�������{���0i19�!n�s�>��c׏��Ta��H�d�E|�K�����A��D}(\�ƽ����Ѯ����8���&�I#�`����>/*a���x�D�CI�#�/B"\�ªxੜݖ�~n����:6��ED�â�Zg��ֶ�iXm&;��|���W󁎑,ˉ �a����aH�?�D2�heC�\������+%���`�Å�1ͨ�{�s�	KB5�={Ǡ^�y~%�ǭ�qƤ�H}?�#)q.�������������]�� K�]�3|���<��^���y^�	6�N��[�g,��ĵk�8��������o�Ut�E<���)Yn��)����|1�9�+������+)�B�f:���ǡO���j9:L�M��5
�n5�̖�^Qri �67�d;��	0��@ܼ����K>)5n�K���::�< ���wJ2^{F=5Y��V�F�P�	�6���P��ɕ�9�Kr1��{�b��ucʦ_9wd�ʪ��#�J��}��sNɗZм�`�d�֟z=��>�|��1���hO����^�ӗE:Rb&S� ��\�"~<��	V�Y��w�W�f��k�*<����릫����6�r�!P��3zA���Cs7�[rk�L� �iNv�Y������?U��E*��'&kC�a戶�X,_y0�٧��hRQ��/9G���UͿ�W��3�x���<[����l�E ���W`�� �&zw�|�Wr��r���_�����,���i4�
���!:&�Sqn:գ�˟�E��nWn���s���
q�9*���ֳ̢���nǖ;�����	�b�x��k��IE�	8�(L`�e�n���Sp�=��A��۷��D#'����y&��@1f��쭯'�F��&W?G�q+��"[�X��%��rɶm�g��W��D����|*�^����H�Ə��\Do��[O=v�?�?�}��֬}�>M�}�V���U��X����^�NkU���hgQ�بZ$R�b�&	afέ{ȴ��.��4vB~C2IZB��=�!jC�K^^�Pt��6�����R9����;�<�ۏbKs8��ͩD�bB��$�$�?��e�j(&K�^W��F���ƏQ����ʵ���,���W&��m�a��ψT��3�X������W§���<������h�@�:ن���z�P��c�0܊��Xܛ���y�����a^���Q�����U%��<�� s��/��v܋�M�OP!�Kḳ�cۥ�j�@�0$c/W(Q�ϋ�%�y��睑Ox��
���n�����b@@�K�Zϴ�c�"N�C6d��8��8��6������ɰ�ۋ<��:��c�O�¡��d�t���c��Ե�G�>l���*y%��b�\���9.�^�� #ͫ�U|�a��0�ea#� i�[. � 7?�����l�jZ��!�#����Z������#���YC��1������)�v#����NݧY����ջjB��'�>�!�"P����G�Wsw�	���6�	��U�v����g�5��'����qf��?��͌�#�0~��O�/�r)�w�k��E����JN���������ދ"��P��i�z!���s�*܊�ϵR�Y"r��UR�T"��Ey�Q�X���_��	AV�ի:D�:ɴ�Cy q���`.�'z#|՗ǲ �� �⟐o��.�`� �M���������>��l�zY6@_G��,^�*��JY ,q|XX;�$��a�-�0*71b��Kh��ӝFA�����euU^h&?�M9���O�c.����mRÂ�̕�O ���w��̏9jL����9�5@I�"	JYd��P_�C1Nl��C�$P2p(��s~�����@��F\�ɜD,0B�C�l	�<�O�g�z�I���e�������<h�� C �H�&��z�����5;A���I�|A�M�Kb��~qF"׊��ÿ�E���/�ǌ{��%N֭��H�Cm**�������:֓yu��-���F��%c�dWin���'����_�E�9[i��>�m��J`F�508�C��<I�����C�\.�[��o�]�h��Z�_��ك1���7t��D���/Ρt��[(e��Zߒ�\�6���vo�챉eٝ��]��fҀP�#�Z�X��ՠ�G��@��Sv ���|��y�����M�z�+���:0�Q��{�y���.2�X��x��)ʛ(_�0�]��n8Բq�^�2N ��N\���Bܻ�@�x?3��W�U(i�+=�>2��.�H^W��[��P�-E�]�}���}�'״�jG�W�n\��0�w���/>�Z"�i��=�^��efeMk\l�b�]-e�f�(i$`/����Q봅�{��z6c� ������V�n'��1f"����(~�+�M��@�,p �,>-w�p-DT�Z����΍U���9��\�|0��|0R	�2���^_^5^��'�;��h����k�,k�q��� O�|rB����>y��`̖uA�P����m��D�/���Φ���U��KJ��h���,����c`�|��q��FI�|�ן��o$Ƚ�7a�6='Z���7��Z\j�Xg< g�y�����H�5�=�@���	,m��"1 -ŮZ�?Q���a
J���4<��S�2_��'�P�<e��˅&�j��FR��\2K�-I�NO������-�2g�e�Uqd(��h�TUew� ��e�j�kN��wŮh���p:�㕃0�-�6�ȖM��(��A������VZؿX��%ր��8YZ��č��-~��33��s�5㿾���A�L�[�l�K��Mc\<��r7���e����W��񵑣���ͷ�'*����$��iߎ��2SsѭH3J��TK�P8��Z�} ��Lt��fس������@ԡ}3����>H8;�s͖��i�z����8�E⌅eG�[��Ab�g��Ƥ)�i�&,Bd��(E?��f�6m�~pŦn�s.g9�����:��#}���2Lp����6�.���~a�>:_����a3�-E> �U$:?�,�N5 ^޽�>�hc8���%��Jy�?n��P\�����X�qO�!�¿��ʙ��ї{'�m��L�SS�O���If����=s��5F5��z<�H���j<@^<��J8��5ؒ=V&S�S�6��#�u����+���jz����M�b�:g���lAZ��	Ge�Z����p���������@,NI�����S��y~&:o�n��L�K!��!X�����nI7��4��<wI5����mЙ~�F�-d�g�w��C+kTID
O-1�^Z�]7��u��<�"�2_;+	NS������FW	��J^�<�g����R�PJ3+�@p�<���ͽ���$X/އѿ���>�
�>0Gŝ�F���4��&6 ��L�V�$[z�q
K�?;M�,��^0!5����ֱ�%��������_����j)ͮ4:�|s���Mr0�.0��S�?x5p ��^��9�|CK�Ԧ���)����9�-�\�汕��&ޢ䥍T�$g5c9v�,9$��6{��
6,v<�at/�5���"��3:�Iz��ro7���>W�aŗ�������a�+
Kg�>t�!����쀨����m�R��N>�s��^�k��Ӵm�ܫ�p��%^<N8U��(�P�M]d}m�
U@#EHƜQ���q&(���J�@R�d�����Xq�G��]D��RW�����]�H�iT<<�h� �&\�Z$M����{^Qڇ/��4��XX>����n��'�7��R����0)��ë����j����4���7�l�d��&ږ�?`������l"
���1Ck�*u����o6'r�?}q�Р�����#[�)�)]~Pd���-������l������eG��c�(&��q���%���q�f��$���<��.��?Ȃ�8e%����DS"��E�q+tO~Jg!i{K5���ʛ��d�"? W�A�F�[��J	�XZ��DY�I^����9�ҙ�E��Nr=;3�����CL$豿�9
2h�>�ݕ"PV4�ZR�i��ܩi�u9T�M��N^���E��?ķ��uq����<�}|h$+�%J����·z��v��sI�4�|}3���.5$�(�GH�1$J��i�[3Nʡ����?��e���Ƈ[������+e��
��3>����G�}��LؤQm85ڝ���2a���!?a����"�Eu}���>[Q����3MMu��q�z;*��DJ�_"6CQ}ڱ������v$�/��y|]�p �ء�vǇ�4�l�z瓮1؏w�rM�v���O��FK��Q`�~l;`Z�(!5�_�;��qrw���7L��F���wܼ��?�R�B�z�x+�̄�<"LU?�N�z�)����A����8#���Яi���D�(Q�<w�(������唿����/��_]�����Q#˧�=��<p�,ㄣ�Nn�0�Kc�V\���1)
r�&�zL��B��T ��Y��!;�s��h��tQ:��Ν�R�L{�)�]���Fc�s}���p�w�Z�J*U�{C�R�X��/ɏw��9fWMo��)�g�h'+�H݁Dre(mL.��3�M��)۹�@#\�~SX݃rf�臟/'��n��K,?5�m���:�%[>èk�t�?�E�c�Fag+f�]�U��|�;0��|�4�1d�-۫8;g -��<���
1�A4�7�7N�`S8I�sn\����TɯT��5B,���K�G���^�����ő2mǫsֈT�4,&���#���UX�%�L"�7��		D(�9G�F����.%h���DL��q	iM�>�hM�|@����`�?y6ҭٻ�(�sE�s�E. U�.���'�I�pn�F_�/E�u5m�-��*r�q,R���޵{�������B~Fc�@H��G���R���k���?���5l{e����]r�-�'۠5*��3���jz1yb9��[�<�T&'=�r�rzV;�X���m�5Hm!!�4ODY�t�τ�����L�����k�j �qM��A�7���01fge�;�#g�-θ�bRz'w�>����"���}O���?����[M���� �� �
(�gFc.�i志g,(a�Lb�4�B�ūUJ��;�J��6��Yk�B�ܔ e��[���Q�gq���ߒГ����� �Ԗ"��g�w˓�.j����K�n�%�΢Rz�@�̘Da��/z�����le��2L�2�>|O�^O;OW�t�N��9�[2)�I0��"�Ϟ�]��`�6$w5��e��+����v�L]��Р���u������eY`cca�$����[0AA�rVt�P͐8�>�`<S�IU## �]�ծ�n'�5V�@�rݮ��TT*l��(��mJn��=�Ks"��� 
���~j��<���T�����f��r%M�Xé �����"6W��Wk�gՕ|k���0��IF�F8��v:���v0{l�. c�{z�W���L�`���NR�;��3?����I*�b����,ۮ�$��@��s⧺��=A�9yD�V]�$����QP
뒚�t�^@�ڃ2��>_6mN"u],���B/>O���A�7�gz'���;�1M�/jj/��/��� ,^�������5�.��(��|�ʎ=t@��!J���'���	[��?�� py.'�o���-�X�Dy���K�le�kY���g�k�o�(����&�^�>������[Z��@�r�$���BI�`��a�Q �|l��yj�J	�/z��	*�d�OQ| ��[�xټ�/ޝ�$�i��F��o("F�*A�k09���\�i��\��D��Ji9^tM���q��4M���>q� ��q�2L�f����;߆4���E�܂wUFg��B�OaV�+ �Ǯ*%#Bm��&�+wO'�;���
�����x.g��sh�7Q��v+�F���[��2Oa���v�c��ge�j���	T�4�,�>�Ҽ�c�O�{2&�8��p�3��Ȝ{��3Z����qBы����QC.�
>�4Lk����$c�7h?}�/��J��Ie�K\��!Y�cb�j�l�y��y�׺Z�&�Ķ�*\������|��B�~���= ع���T���!����Ι%-:�ɩ�1�����A4đ�����fv��,�xNƷe%c���"8t�>�)��:s�%�9:)!���H���X�]�ŀ'��g�s�|�J�ş���44�$�;�rcs>�hR6��'�������I�A�����.+�ǋ#I���	]��l���jFs���]gWQE0&J;���S �?����^6&$w�۳������	9@d��\�?�*�a!t��؅��M<�az3U8�?��?D)� �֐�����om�v�XW���d�h�K�/g.te|2+�#�D������D��ãt㷠�{���O�-��@��a�Ѐ�`����рH(1���k]|��^�J�K९� ~{r��R��vp��Q���=�'�����!��k�1��X���Z�U�m������jS �����S���Ѳ�k�%��Uu#��)a��Ę�,��N,��6f�l��⟴�4�c�1��G�����lq�N�4;���$띗�K��U	PX`�&��v%G����T�Gp������쮛��\�(��m?~���{Q��j�ٍ%��(�C�����ԋ^�&5���F���Yā��
�*�靔`�H�?���5�Cȶ퓢C�
�,@�b)��*�]T㑝�3�6#o�_.�!�:��_�.�Ҍ��uѠ�N�Ǭ�sV6�'���H���Ԙ��b�N��^,)��m�rP�f�X5�L�P�?�M(����E��a@��]L��jK6e�6���'�i�$����� ��ġ�K�,��e�tȍ�3�<B���Z+���Q(z�J�tt=���f!��j�n*wG�yFH� ��FG��3X�ǌhN���# ��\�E�N��� ������n����d�JAW�r��|����W�͸HT�?�9^���9��6���W��T3���@E֯B;���+} <�������3�"\
y� �3f����W)�Ydd�>��	��;!gK۬�����d<km��S�VĉA��}W�	<t	��<��)�ժ�4)Kb�8��&/⛓n���#���z�2��*��e��Iqʹ����Z4K]��c��u�����c��{Љ] s�(�� ��v��+�M>))��H� �i����ͥ����4=�3�!�C�{F56'7��+@X��M���\X�ܱ��7�D2�"�T�s>N�a�6��_rI-�2���Օ��L���|�p-%C)�=oRvu\˄_W����0��:����b1}�������ה�B��"�M[:��
�8��=�7�/V�c6�㩐��e ��f"+K��U�X��Y�{<�Kb����:�h}s?K����.�}
��W�OXQd��D���J�&����ໆ���썘sh \�8B���)��$/^�H{��=�� ���Jy"�x�]s��<�0�e�/�v��BR���o�-3�Y��2EU�ʘ��z����\ĕl�.�f� X3l0�]v;�>��C2�w6=�//� ŎN��o��7S��Ƀ�I���=Y�.���#�F�x���W�2`�y6j����`�L�RFh�f���0$*EN��[���;kV&�D(`�jo�?�q������Lm���Zj�R�����r>�#c�6eLF�D>�zu� ~B8��Sd(i70Q��M��?���\�F�g�������jbKX���'i	M21��BB�5�s1 0���(���6+�xf_��%M<�Ͱdܗ۲w����E >��@~�]\�v �� ���/�	���O&NA{�BC\.�`�T�� � �t��Ƚ��J���`�p�4K$��fC��k�R���?4-ʦQ|
U}�~�H	�ь�ž�t��5p����%�
-�7�xw���~���P3�����?ǒ�{��͝U�.�mE�����f2%��*bk�;[���ZT���zW%M�!�ǡ�Ώd(G�#t���ٹ �  ��E$ͧ�؞�,��l��I�yO�Yds'�%�wqǆ���F�f�u�=m�Z$BO�[Vzl ��<"��p��^�9�q�0T�X!���֘��UC�;v'V�6��ȞS7����<�����K|��M���|~�'ꆁ�L�C|.��;�s8���|�u�6�䯟��a��_�^��+�U��orv/��';Q�O!��?�5;�k$��0tN���͏eÎ���.�T���4@�K��^��y��n��r�/��m�\�X�#��&�E<l�@Θ%�Kf��`	ʮ�Zx���tT�dQ?�{ ��Nj��z;pO��x�_蠳?�C�د�	�)Ӳ���3�	�ذ򨹃V�~�<ޱJ���PV�2� ��(f�"V�N߃�C/&���S���5V<ۑtS�Y��.-�Yr�� A�4���P��8�=9���g��e$�ٱ�.�[a^'r="@ӿ�[��@;�'�sǻ�,S��ѕ0��/�((�S��h��\X�txQ��,�e����@kI���5��j$ #(C�v�W��'Kn�'o����-�LW�i;ګ��@k]ќ�rò��d�ޙ��� g�0�V l:@��u�.�E���j��t}�a�`���VEN�Z��*F���v��-���n����k[��G���أ����1����]`�}�H�sz�VfZ�:���B�'l�:0y�t�����X��f��'P]��S���{�`4�b���ŀ{Qj�k3����l!�	�I�<�e�o�3`r6���2�|�;A|�/��╟8��MDA�j��Nd(9S)��S-�w���`/X��xF�j��p���T�_|Ʈ۸|�h�䖖ǹ����/XbG�_'�%L/vgÝ����<�R�~[�F1/�C���� �TR��s}�QT�_��J���juY��G��ٔ'�%L#ZG�'���	�����^cd�D|���V�R\b��1�6���F���&����[+�ʭ�h������ˋ�z�zχ�a3H�#B��&���j.� b�]~0�[w�/g��O��Cq'Y)��*^�e��P���{��Ē �RD��Fs� ��s�bT*�N��1�uCenc�ŝ�ͬ�%`��U��FPʮN�����w��$�ʅ	B;�"�e�څ�Z��ۆC+�rq��+�\��%6�)w�����7fr�&z�.wˎѝ��7$p1g�� %te��.J�B���f#�����s�s,d���X����-XXi|�E�)ab�K'{�9o��aS5�SA����WC����<a4���C�����z����nY]9�'��⌥���%�z@�����
��P�*Y�~任�B^��H�$L #2#	Vb�o��"�5�NT�K�y3�Y
���sg�����k�2?�7�n����f�<ȓq�ݪ&����?�����b���^O��=!5�롫�����s�,�����/����}9�wJ)`�Ʊ�Q��;^��L'pV��HŲ�1�[�x�E'D�pD]ʞ�A<G� ~��o�p��:�I),��Ā7�^R��K�鱒눅gx!�\���+�@���1��g�����ƹ�i�?�hdc�[��uvf��e��pW}v�m���oY��rh1e�oX<jg]Ήt_�X�9g�S1���R�bpT��xg6C�n�%)�^�l��.~�V0�[i9֩ڗH���jG_��ݱ�H���k���_��R�����@�.��TuK�ϫv�t�I���p��(AH7�n%�7fȈ�âG$3>o�X�yi�al���aX���� ��PP�����K���L�L�b'r������P��s��3\V�yB��+���:S��Pg`���L�48�+Uz4���<�m�+匸����җ����������M�u*ݕck�9�T�����45ۺQвt�oؿ5����ڝv:KB�/
(� H	�����2ʷ���5�&���~<��7w�/�<Y�G5@S�AOtq�'��[�)�W�yґ5�H��,C�Uq�i3�����اQm,��pFcpW:$�8���U8�EZ`G��]T|kɳ_���{IY?6������ȡ{����C\�U�3J$�{�c�5M�/ܞŤ�Ɗ�a�a��F��qFz���[�����'�c�N�o���]�d��$�	�j�$`�N�?�X�e���{liyc�9������5�;����#/}���;{H�Z�Jk!���} ?0Rc�"�E�|�G���b��kl�o�������s�^`�ELU��j����S��l?dk�����~�{��1��P��e���m��:4����&l��������@�1{�n���Q�o5Z�=���5<�Z����xL��n�B�����rUD�;�/�>ZD��UЕlى��ѿ+�,5��`��N��"��@���t@�G|y���L�ݵ����٢I��Oc[K����W"��Ӣ��4
�3D�7�+��K��G=�W����`G�p���E:�����{��T-`�-��3[rE�[c�8)i8lMU�%����G�܄gx��RY4�G	��������5�znVpM�z$���l�9LI��65 ۳�= ��Z�_���g��\9�=��d�����L���%���ת��r���w��х!Pwᚓ�˄.�~��T�i�FU[���r��O��S����#yU�:������eX�E֋���O��/a�m޼iٲ�S]A��"�O�)����� ���q.]��JQGa��6�
�e�p��| �?�n��.b��UU�����|�e��"���Ci��A�Rb�H+>")�(zvP���ibs�n��2
>w���x�R� �Y�Cie�z\�d8Q�D)w��%�B2?�帿���W��NwЋ��_'Op�D���ۥLaǟS�X�ڰ��̫������`�g"DG������u�׸����;�[�,1�������_���Z�j�C�ġe��DlHg��)�	��~��x����U-2r�J��?w����գ��*�SE�`�T�M{)v0?�Z����-�D���S�j?�Ao_�^�2)����6#��sگ���$�03粒�g%���&�d�nG��0]�g��bO*h�VyA���d�U��q1_iK��9Z}����(���?�b�ɯ.7����2FB�-����Y>ǨOaPZF���ilKʵ���RT���WS�m�N���=<����z�R��XeF��dWV�b��^���{���M֦������=)��J�c�j�x���s�Mv*x��
�ˣ�fԳ3��w��i�5���I#�A4܁r���@��b*��e) �F�)�M�l�4F���g��s��o��ưV�fS�iO4��2��S(����8�y�W��sWݾ�"�i��p(��!����%|]㵙�^H�Oy���AQHPD+N�2�KK6<�x�XU+ɫ7ړ@�h�F�h��lT@�I���7�!f���`��#������bpx��E�M��3_��s��hL��M������KKME:kKP��E|k�V�FŬV�Y|�Y�4`n��ERi+�|yp�>V�/��E�i�s�>��+/������͙vE�2���,m]d�gU�f}�t>MQ���aP��K�[Z"�����KB��˔�2Շ���W<S��ޭjf��%YE�2�c��� �x
���Q#:<�d����c�'���l\��վ��n{˼�-Y(T��΃�+�*��+j� a:��~wA 
���6�; �j�Z����9��d�q�Y ��/A�2���b�,�|��g�u���3j����xo��<g][K��t4G[���D�݂͎�x[=;�=V��i�R�����%d�s-����Sv1F�/�s+T���0(������!%��k�з*��pn@�r�{��5wz�	����>�?wN4��<}�8�{v�eJ�M
�g�Y�*	`Rx�7�Y&r�
[���{�����h!��?��h,������L	��ũmZ�C���?��&
d��$ #��L�2*��;�z�D�r����IЊ3�g�@Qc� �l�ʑ���p���n� �X�e�!΄���3B���I���1la�\������f\1����U�[���k,��Ӝx
L��V����礀���Li��q+Х��n��,�����ZF��S�f��y����~~i�����:;����c<�����;��r���>��)#P�����0h����4���h�q�H9��aHx���q�1����,�g8�?v��*���ם�lj�	�T�N� �N!��'h�ͩ�؝B#��Զv�����(:E�9i��[��5a$�z�O�%bA���R� ��`Sr��\S�0�846+��4%~7����	eE	&���B�H\y܂:о9��M׏̸~���mB��Y^�e����X�r�����3|��6J���
o�[���%}�S��;&�#3���q%Y����j%��F+�^iv�?ra�W�j���v��A�jYb�Y�d���0I��w=1`����`������v<Qn�8p
�3 pm!~&<�[eZi�����C^�����[�"��]�\����%���V�I)��m�ŋ,�rj�9Z2]0D��\L�i&u���&�HiFM�J(��� ��)�6��Mq���L�?�ׯ��0�jn�/T�v$^2����[��HU�9GG���~.��� �g��OR��%����oU�P�TL�L-&��q�y�>��<�lA����Fb�����*X��޿mX���3����7:w�t�x���VxJ��n�r/bmW$��(���Բt�vGec1щ�)�'��)��D�9,\bM��<a�>�l+1��|��\>я2�-��1Dc�݌�)/��Y[�=7�+��̿B7>�@��$*�kȷ��LX�"m�Y,x��W��l��dL�,���g���I�DL�p3��|g��Hk������	��>�
~214D��0UM �C�+�߈�,J��5����#���*�x�[�8
�J�y��K���%YP�3�g�	u��@�K(*�WM��� ��
���	U���4b�΀+����|������O/�7M�,2跰��]q!N�2�Gc`>PH�89�;�u�e@+��7h_j�����H��x�w
k!"~���d*f\1��}���U"��&*9�d�{�)jr��sm��6�+"���a��ƫ_f0��^B-3M��d��?a�=ɖKmy4;�������:ܺF�b�ZV�*2����	�z�9Kc��#�T<�R�1��ڍ�����#�C�SqGM�����Iؼ�&��[}9��n��}�b��7�Wo�*��B{B�h��d��o��5n}�sp,�_	���T��7�|S�� N�w�!9|�{�ۑc���Vn>�<�����k�h�0���o�y~�b��_�H ��OO={Q���e�gQ�;�&eh3��M'��LI�
�|����[su;���}���d�M�O�+���'.�
�4~e�쇑�ӹ��/�7:p%�e�����*�nh$ߡ���Z}�^V��&/4,�l���_�^�b�'RG�{�K1������H��?�[����$^�U�/�k�R
bV��|�F�d/�0�����S�[�@x% f�v;F6��>��%��T�
:�ë��Ј��(ε�k�>��8!�S�'��ϢQ��#�y�O#��Յ�u�f%�&�\�Q�<$⟥����\����z��,�J��e���mdj�q�;l��W������r4�h��ga�U�=��D#܃gQ�哩5V�ވy���^�ӍQ<�Ͱ�̾e[4[� ������p��i�{�|�?������Q�|�K< C7��8��B���o:�Y=��-��/��u���0S�JɊ.�A��^�5�WJ���iN�@��-����a?g.�I���� r{�Hɾ{^:�㕙q#k��<FC�f���<�r߶�#��IT���$����Q����C>�0�a:�tYA�*���Lr�8���B���^�ˍ�y�ȹ�v�K��dH�e�Ь��f]o�x��&� /�$5izEUL9D�S�Nm�_��8�y H�f���!p�o�xs!��rA��A�$�?��YG�*�K�M�T8$�0�<+���d�,�O��ޞ���g�D�ApED���,�)�R�G���5��6�x'X�
��p<�X	|��jG���BQ�� ��G��W����MG^��7��~1��Gy�g3K���v1�[�����Τ0�PkX&���\��&3O�܌�d �xW�+^*�,�}��d�4,�A�bjrI%'���ś�h]P�4�ծ.�;�񧢋�=8,w�mF��3la�N�=���i35�M����"�q:v�9~J���(��/�RA����@-���-}���t�>/�$A)��Z�-u��L2��a�]7����6���uj�O$v��1FW/��C/���ݝ?{�Q��G��-��9����Q�����\�'��(pmɾ�H�2������gʽ���O�Yx�!�:��b�"tx�p(�L� ���V���&�6DY����3�O��&�	+�|󆄝�f�#��l)�t�9P��*�Ičt!��W��}����,L2_�_���j|`8���\�ս��(�!�`5^�&S�<�+]��2jOѶ����/��O92�Q�O躺��E��]/ف��{4�Dr��Gu�9.f�;��&��\�ɤ*P�W��6c �ԧ'�p����@jX��Gsޅ	*�d�S�:���]C���۾�LCk�V�{*���9�?�g���ɧ�་�u
�0	^)\���[�H4����'�	Æ����0������ޭX;H�Ki�c�TS౺-P%��_�wA~Ǻ/�L�_���qS��+%�r�RW���q6����9nn��d��6�϶��ayGK�ka��Eҳ��1MΫ"��-��}����G�c�p9&H<�AFY_x����V�xl��;�
'�{ �X��L���'�]�`�$V7!���L��+^���;j2��1*3!7o�+�I%���>�(���pp��łD}�~8���޷H��"n�5U��(}M���Y/+��W�)쟴dv4��{$�0���JDO]�F��N�Zd���ϴ���}X�\''�t��A_��{��c�/��X��D	�U���=|��`rz0��t����Tޅ��=�%U���QM7<�+s1z�#Z�a�!@���\��B����!�?4�y#��]�O��i����|C��!��k�g{���X�r���M@�{h�)������ꋪ�P<�I���I��,��>���^M�^�t#��S��c��5/� F����եV�j�c�Ht?�<B^�`T��o��'�x��K�D_�2�R�Jl�5�F�*ƫ��<~����	��v��*	����Y�{|Y%�ō�G2=@(TV��X���?g�����hY�9.�b�
�}��l�g��km��B�&~��PvLs�B�~>���P$�^�R[�}q�Kk����F��<}�8����Q������ٌ�����
O�	�sCLIG��d���1�k�}���>�-d�,x|
�������%4O�QZ�`�OP����L��w�'��ja_�N�%:YJ��g~+�#��D����R���)��۩H��ٰ����O�PU�Ջ�b�m4*esCr��c���*��p�� G��8�c��ĕ�������@S�׌�z3�?�?�Y��cb�����6�"*r`a��sRǮ��R�����I �t��U���	��w`x��'B,�HO�� n%=��m},�ir�|�l��[��8���G-<O�.@�/�3w���E-g>�p����*�����s~���˕���
&��#�qZ�|�a��)}���9~�/�2R�����[���K�J�=ZCs��Yrݡ��<�H��_M�z�ͱYR�&���U���ۄ�a����d�U�W���5��%�D��lHۑ�T�Ϸ��t�����'���'��F�r��Qx7�+�Z�-�C����>�����'������!��:��*�y;��x�!��:����a�{�4��;���V�'e�L�W�1�`XE55����x\����6J�.&���g��4+l�f�#�{���'o�rߝ{�W�9F�wF�I<!�N�� �*��+�Skw�`���4d��~�����RH��q�!��"��k��m#�p��ѱ	`H��N.=��xm>͵Fb8���Sv;�a�VJ��j�����(d�����wudܸ�p�tÓ�뽌{G?ߡ��	Ď�LV#�����;�M�@��?����,�,��R����SaS�Q[����yf��>��.� /����^��SҎ@6��M�ch�*�nMjEi�H���q�����'o�yC����d��c8��FϚ\7W�2�b�͖��,;t�1hJ�����W釼<�E�eQ@��շ�7��\���,z�!�TVq22z�Ե�v����X+^|�O�*�Bt -
8d)����y ���a(B�D}8�q�jd0�v#�kg��`n	�m����Ȣ�
9��~�y�|ܣCG� J�=��T��A��']���M��G�i��#�Y''�T	���ّ����/��DNEC���W�|�q��˕3��Tǅ�9o�8�,�*\�aN��~��[�n+�$Y�dc��BQ��� ��c� ͆�ޚ�t�4er�Zi�Sܱ��D��2C�J���u�Nc�����˷c��VҶ��J&!bagi�n ��)v�Bӊ^b���Ճ<�0�v�TBɕ�3j�Z�jh�'aOH`}^c3�M���8����g�b73�Ϊ�W"D�ǹZMDz,b��z��J�-�´M�a����Hp������q�爐��g!�1���h�(��Kǔ�DƃEN\]��h��.�3�Zk�n=x��,/��������>a1ܚ0�;�)}���^0��|�/��|b�%$~;�	P��p��ެ�3�m����_E5�D@^�c�ܻؓ���v�fE�U����㪠�T4A�`�\�p9���v�K�0��«�ͅ�?�H���"V��
C�����\��<�$�Ϗ��k��+���"x	F}-}�& ��lߨAJ�'U�C���H�f�p2�>ɰ]'˜ù:�Qr\�N�"���`]z���%��1Hbg2�;c�A��������u=��VLQ���'��b���(H2j-�5��L�N_���XvS��ȫx��2�hqM9�c�/z��:��)���u#[#WC��M�R���xE��1*�<�����ա3R� >D0�j�o��+��kl`3�)�_��Д�k�L��nϚ΂4o02�+�ֆ����#���I�w���
TP�㬚Er";�2i��K׸Y��F�b{w�=e�����65�W���I��}�o��u�D?t���c.��fϴ�e�\V�:�
?��й.��" �oG&@�C�ē���-�5�L��揻y��Sy^´K	�D����[��DGH^��s�A�<�S������r<���q�t�����rG�1)�����☪C��ﬡ�6L��b��A}�y�$���_�V���Q����.��k ����N(�r}С$6���e�����bm�(B�Q�0!�!>n����߬q;��ZG+n�ӉIK0��^�����nZ�Ĵ�$[L�LOո�s��2Y���Z�2�u?	C����ט�	�It�?�dP�l�L�����o���������`"�$�s���u/ѵHn�Q}��������%W�F������p%�4�d�
X���V����e�MJcR, R'��/>��R�4��p�ŋȺ(���x4�#��Q�h�Gzg!Q����0g��Y�d�	9�b������ҁ�ln4����V!�dn���c@�`[�f�uI�����s�@�Q���Lٸ��(a�@o�u�c��vB�@�@-`���%��"K7�я�����5z��q���F>��oBٓ䵹�4 2���nB�k@�z'�K�n���b�����;dLp�ڊ��#�7�n�6��2-�8`�#V�%�SS��3O��/�	��2��5YP����:|��w�[#����Ր�n�Z���őGPg�-�
<�If�'���yƒ�O��~����+o�rc���"/M�)�Lk�^YA�M��LL���sYJR��Ļ?R�<}:w�xG �iH0	)� ���`�_�^gY�LH~	Kw�,����!��VW���H�������G4[��3�֏<B�I�޴n p�u�Z��'N�3Fa'�Sn������uT��`�y�NjV[K��C�,-'�G��M|Ó�U������m��\A�NPl7���0y&�҆��9c�sP\z���H`e��V�?���A���<���{�$#d�{�t���r��J��4�����\:��,i5��W�<�:	�2J69&6%��1�saO^�x�5�y����������F<�x�p�[M�X�&�&#�{��S�9
.Lx�F��p�I%�0@]��9�Aˣa�)��8�%�H[|�'J�����*2ڙN^e2�R+jTHO�u���pI	�Ks�ՊRHu�@o�d+<�,f��gp^��s|K�#kb�Ց`�e�q�C�ߞ������y�Nf��c!}��$�WQr����[AO@]sܺw��w2L�r)�Y��g��ł>!�@]��$II��֯x�pd|x����!���|%j翆�,H9.����	( 4K8X/�Sg5�׈\y$2���Pڪ(���j ڦ�M�s�*V�Zͱ���|B!�g��V|���3�81D�K��w[�?!z�lm���.ψmX��j � ��<������_�O\�?��Yc�l���P<�����nD;���������C����������6z�{۱dh ����iڔ�XR�{�_���}�0�谸��E�˕�V�Ƣ�.��+��p�6栾�bF��cW�S�@�N���R㴳L�s#��D��cn��s/p/����4\�s�l. ?�Cn��OJK��X�ļ�_â��]�*a]�?��iv��'�Md_�����ƵrI��Yj�&��^EE[����j��=��W�o��Ѧ"s{V�}>V�g4�ِ���`�d�,Ԧg��5-=���U���+�?�2p�,
��2�������6�Ө���vh����+��Y���f�+��mܰm�7�7鞃���j��Ce�����F��k��?��#�!��g�ɷ�ܼ���AwR[�>B�\\�(���)�OZ"���I�n�8�5d!�����y��j��[֌=��I�rpjC<;~ѥ6�/�f��=J��.�N��� (e�)�d�M����Y B%~L�K<�r���>F�q�V�)]�A�F̟��xЅa�����xUJp��P��jr�u"�
h�r��$觞]��͕���
�Ae��Q�1f�B���@�¤�v!�����s���2>+]�m�bP�T�W,`&Fv>:����D��I �rl�ml��O�0�݋o�i	4k"X5Z:�,��ڠ�Xzf�:�k���9�]O6����P��jI�N$c-��X7�D��]�Q � l��9�K��̥,j�F0%�`O����ϩ�g&bB���\>��#��HQ�e]������T��Cr��0��z�_����1士�EL5Q��u��I���ؼ��hy|y[��t��0�}E�h�Ҟ���ݜ�7YhLY�b�>-3�<ܘvI�L�e���rr����F����>L@�yjF�`��Զ�5�j�I?j��}�ԕ0k��I��&d�<���@�5	$�-_�X���hM�%�v��c���{X�b`��Y�F=r<��= ܨC�!�Z�������+�K�R���m�<�6Fh���g�U��l�=�NrDKO�����`��1Q �N�ɱ�^�\A��+ܤ4�F�����']h��TA᜽�_��I�z���q��}\b����锁K��"g
nUiL^|���19�`��H�p1ִ�Mt4
3��y=��Q�R�`�@
��F�5O4���֭�O��m�w��-Ԭٵ��6�F�Q�CU-F�z�X����8�z��V��x8u5�v���\ٱ0l��ֵ�<��3c$p�윭��,�I��+a�C����*	�	mK�'��*���zk��C�^����[����7x�k��B1�^t d��5QǒQ;vB4א�9k�o�A�M:�rm?�э,9ܾZ�f��j]�u�T���U�]f'J�XtN��ؒ�}��A��e�դG{�����&��a:����v�y�wY򐘣>G�RŀV�}v�M}�B)����:@��g������M�E��м������*0xC�3Fo��M׭s���*�l�e����I���b;Ftt�kNǆi�U�x�:ꂮ��%�)�~c$�g���]v��:��DO�g���:�1f��w��o
	U�.8 ��8�)���(-;�� �G�T�86�_E4Fr�B�������Q�QJe�K�-�(h���=|���H�d�[U������}X���b>n�w�wS�PAL4I4�g��RX��������;.�ʚdCj{��ϋj-߶N�i��fn^����$�˟�*�u�ͿD,<������[�����K�!�S"����"�<�m��� ?�����_�v��]a����M{�\�aU�A?M.`��|�v��O�]�'�'�s�^�� ~+����.��g%G�+�-d���S�h!�F�{���rn.:�� �T��<��<N�5�ur죀ږ$Ģ
xg'⃉���W�]����艚�U���U'����͍#2�gHN5Tى�������3X����=0/�k��mF]I���x\�S�M�}ЀǶ��;����_[�c2������Y��k�G�Gv�/�L�I07?+S�=1����X��oI/��c1��f��H�\���C=$l8�z���$#��0�<���h��bz�Q�a�-XVD=ƾ�]�4�C�8#��`�������P��;��ڳ���zH	�8!J�e��u�	�̖�O(��Bv�����l�6��an^��!��?�d�:oU��H>���Q<��-6Q�0Ao�0��,3�.�!.��`��r�7��z������&͗!�mK�V�q:Rj\8���q�*�2����R�2�"!���9s��Ah������4L�(��ȾǗ�u�k�����[����D�]�r�II���>���Kp�>�MQ�pD]��ȅ�B٫�y��Z=�v��� ؎���E��G��������h����7W���Q!V���ctB�̑:���ov,H��Z��z�$8�$Տ~t�'�/�)6+���;\�$E4՘�󖗼�SYn�����v]�-�z�LWO�=!��>�g���o1������	�:3�[�${�V�s�o=_z��O#����e�{׵���uJZ�u.]���0 m�g�]	s�m����F�jC{v ~����+=9�P���cu��8^��
��@̀���Qf�ޤ�����H�ʴ��k��:&?�[�[�w�P�k���M�o�֮L"b��������V�=��P�x���������FWa�Mrj�a��@��x���Ρj
~CP�ijτo��� �w6����E�?Ɨ1��Sr�d@��s'E��zĥ,y�ԓo.	 �g#C6��G�٢Q�EkG�8���tr�|����2q��cK� `;�=�Ӽ�����$#�Km���;,����&�Ś2�}p&�oE�����C�FT>���Y?֥�X}��3YX6ɡ`!�@�L�rb+{���U`�l�#<��.r+�B���(�#���4u7����!B|�&h�~����~;�ad�#���;%rfԭ�7e+���L��@^j=,�́�AD�u��ƿ'ܜZ�7 )��R��j<N�A�5)K���0✄D_H�,����$�+�,eз�rO\+��9/��B�R����O��-ﻰ|)S��� ��'A�tmԳ"n$lE�4��FJ�Ñ�Vd�q2�
�-g�&���Og0	>�jYQ`�5Uc�b �E%N �aƏ��w�A^����^����B~�џ&l�h���NEF��i���{�fq�J�Gw<�/[�<�"�� ��p6����3�A�`��VS�c���=�}kׄMD;�8�w�s&+�1#��G�^�����'��Ei�D�w���,6@�:8�|�<��L����lܖ�"�b���^�E�b��Y�� Rn��Gk-�$v����҈�EMp�i��z��O75$�q�q��}��T<�*�P����oO`�0U[E /�L���QT�F��Ic1OET4`���aXV��_O�"AJ~�*ooV�6gŊ��47>&�b��BP>i���=
Y���Y�����Q���93���ڎ�� ��bi?S#J+jT~����P"�� �D8Xx+��Kp��V����?�ճ\��ʢؒ�`�*ʻґw��QZm����ʩ�e�ΠHG!����CT )p�D26
T�:�~�Ve���d������?]x�y2��:�V� %����	������}�a�n���Dx9|�a�h�M�P�g�6�0%";� ��#�0�(f�#�W����M#�d�K��әҖ���dJbtV���<�0���ϘY����2�Q��̙��Ф�
�;��k�aߤ�&�P�X&�8�,�C���뽯�l��<��GjjP���̍���:d���y���5W�xYQd�j�Ao��˽F�d�f�모h���-VhEtoKi���B�BX��D��W,j���O��&paְ�#Ob�S8���V�!w�����V��6���f��� 1��?FT8S�F8�=l�,�؏��Hd�,�F���iQ��0�"{����>m� ��f�U!����Zx*\?��h��J�+��|FJƀeo�]���+�C�*\T�%4�bE@�R��&j�l B�L�VM� �=鄚f���5����^���j�yd��/Ϸ�[D+��7l͛ƅC��mn�p��*x���i��8BA�
:���5r��eN�,����t)]]�%���k:Z�� h�dhC�	X���4�F�,h���ɩN�xkM��v��h��H��i?�s���+�L��VS�OJ���X��ܜ��z��.����|�R~�7�WV�����)�6ms�G���8����ѽ�l��<i�S���V�7@���c���Ձ��a�oJb�xKmK�)P�u�ǈg�5	�*�O|���(�2.S�<�q�Q��J�u�\76s�Rފ>5�u�0A�� �h�>����]���w�Q���'��է���$Y8���lk��t�6)Pr"_����c��XPb���C��<�'Be���P%$�<	Rj�!9��K:H���%�A]l}��{W%SSxz�� �X����Țm5;sq�&b��={�P�\���гR����)X�Dys.A辥�VĹ���b)���R`hw��;h��Q�#|�S���b��:��lU�KP��>;�]�zs�į}�M8����-m�"�Pʜ�=S�������jw�_���S��BFf��ے%7���
f\��J�˚ڝ+%ə��;Lv������5�_,�����>bz�I�rN�����7X�2���m�ܛJ��얾�����hky�f����5�S_��+c^��＾���5���[q]J�ϲ�59�
 ��ɠ���!h˲��f�/|>��J��,ɱXG?b�D�t��7��/O3�R�����RV�P�_a�)�W���9*�Br���R�����J��f�!.��Q�Q�w���w����M�[1Ĝ#���L�Wн[p��B�R�/S0���*I�����/&4����P��;r��+��R�B�:Ջ����]���=���b&P޾�cNĥ���/����߃��
I�V��`	�>�?=��-`�"�X'y��o����K��Bېzk��!F�MY�ѷM�F�c�S���e�B^;=qQ��&ϒ�۞�|�w���R�cX�υ�7胬������1�Ta'NʪG�YzW�7��˺Zr�����aK��e�����Z6��.��;�s��9"���2{22����t������pM1ԭt\⛮~3����;i�l�B�uEvݝ����V���4��_&d��eNЗ�R;�Fq�a�7�3�w�'}"�͹� ��s�~�7���
O��	;:�].��U��+�mb��b�	���Z5矻�ip{�LJ
���k��� ��˹��*�z%��42��iK�رi�:4��1�ʗ*U��Hw�ł��<	9��љ�͂�0�o�V�ky�\��2�j!ԩ��e�_�Ț�������<��5�;/�f�Yb)n"~���fc+�:\H�4��m��o��
�/)��`�@Ƈ{��S�a����T��U�0J�;/zY���o#����2 j��Gc�A�Ǯ�����G[�{��f��AՑ�R詖|V��^�
7���ԡh�%d���n�]M���R�n5VdA�_N�k���cdE�I��E���ٙ}z��k�͓��(D�*;���/֎�W�G�ܡD��E��?��]���� �����wL����\�VD�P2���=�����,	X�%�}��B��A6eymп)"��2�pD-����������~�w<T8Ӕ#��	Ɲ<���&X_�'mz
Wf�`M��.Mˡ��zmhaHm��-Lך
]������H���,��^��ɚ�����y­f]��JhJ�cS�����a&�Ƒz|�=h���_o��U�2͕xm�{d/�������K0	���(ƏG�;�+����@�+�6��֗[�Nvv�)n��E�S�מ��׃ogxx,U�Q�$(��G���a���zv�Cf��A`���z���F��@B/�K��)W�І����7�+��/���ͻR��edBye�\��(��њ`�n�q,*����J��?Y�2K|�3�95���(N���\R�pŔ&|��~�N�I��O'��OR�Yh� %`����D7X3xgE��!���I�s����J���m�5'����[`-z0�U��ĕ$��T�����͐w�`/��U$]
w���i���14X�Ū����û�Ǽc��_f�� iHQ�dr�I�~m�q�1�U��"�o��$xW��]�i~ ~���} �����r��ZК�-,[�Q������Aύ�.�n��
�޶^���'"x��9A�/��Tw�T�b�(��E`�vAD	�\�����I�b�n#J� ���ب��`���҄��Z}��b����W*T�x�P�8�Έ���u$�����]M2�O���ӥyb)�a2J��J�#��@��C=�{ 'VR-W�* [+˟7f6XK^��e��L����������%����<�:$��#v�@@@9�d�D�$] �	ʺ���?�KE�������w����^���|�Ϯ	���J�������Ba�����)���)I/'90fo�u�C�9�p�"�{�?jɆ6uxO�	����\3��?��_}#&0:��]5�=�EA�eH����D�p��v�)��o�!�8����+���\�,�v��u��m�ePޓ�K�W�O�&Bm��f�\^rb�P��ƚ'�MZ��{�8�eL��sP������$#�� ������Dȴ4��>�~���Ƙ��w��آ����� |�|6'o��,X�h;`ѯ+���8-P���_;��M2T���bs�Ю$�$ӭklP�}"���2͒�f#qx�����%��d�7��7��K��(���79�>x�o���_f��&,^E��z������^3�� �,ܒԲ�A�ڲ̥r$��Du�̩?�x����a���f�rmznJqѹ./�=��i-�Q ��J�B
��/ŝ��op1{�	mL�ap�D���� т3RH?���\k����u���X��>?VWP߆T�)�	���|ٶ9
>��W�}�1�ɻ�#�X�櫳�%��d
'|���{$��cՈ��:�ɯNGf�"����ح���Yb\o��i -�{@���ݲx
�y�X3�J]�]�G��lC�@)�0�!ن�u��x���w#(�\��W�#��+_�e/Ź7Xd��u�c��,�{<�4ׄ.M���ڝ��ה�1h�w��Fp���q�vh�20v��ݯ�5�X�g��L�Ad��]hR�E��!M^�x��(���ѳ 0"U�q��{'�>����N�ۤ���r-�A���_Ƃ�׶�����.��b��S;�W��?��쫕*���|��Y{{p��4Śv��S�;�BRW5S?���K�gs�T���f8�x�`�j�k ����c0<�0�7뵶J�o�3�u�^�A���Ⱦ�`K/���*�ڛ_���7�"�L����M���<�q���d�v,�$w�x��yh12e�q_�?nN�V�X������Z
��c�R#��dg�ő��9E���v ���^0��DO��~҄t²
x�����-ɻ�0)�vZ�����$�*G�V@�\d�6Z|h�1Q��_�ǉ)C���fwQ�x���0`�{��AX�Ȫ{����A]�E�	�<����d�vD�1��[h�ǧM�6� l���֣Nh��>���k�b\�P��������ۇ5��A�鮣�y�ա\�ġ��zI
.gZ���:�{�q�nU�x��
Q�V�uW�Q���Lq�Ӑ�C��Qr���W�j��Ӿ	���sd���q��[ga� ���=ܨT՗s�t]��=z�$�_�/�.IU��`M`����cR�M�84�	��9��.�Չ�A ���;��Q�\Ȑ�.dr?X��?��;H�����N˩�A:��&R��3�Lj��W�#t�y�M͌A�� &$2��^��O�!�Dβ��"k	��<���`�9)֮���_'i�Jl��xQH���yc뱿�\�(	%H����'ު�#��Y�L���b2(`�%�!ϭ��(���'c$���.U��ڔ�u#v�H��{�4���:�*ں���E�_/����α❅[`�)2V;��&�'�B+̙P��g\�u�r[��I�ь�'�����R�z)Y!^vl���&ۣ��o�`����V��+�cY-��a����J)�GX#{�	�R����ˑg�+
�Ҫ.<�t�ɀ��Q��g��L7 LL�S�h� �kj,���첐E��ND�ioz:�c���A�h"~zD\x�����'�`:-t�G9�դ����k�Dy�O����h$���6?#��x��S�R8Y�[���:�5��r���: ��������3ɴ�x�@W��!+-�u3P��	�º����i�7��5���O��\���z��j�3�n�W�=��r�+�E$�{��̔,�����K!�<�q��Y�_3��*����D[[��]�!���h����<�j���7)�?���(UD$9/�����R��lj ����K}D�E�� qfq�*ݤ�e(˦�p��죌�e����bҍ��޲�K�Q��y5饐<��]}�U�W)��N��9�{"n�ĸr�z.����@�e|e!��-��&�4�Mw�f2m���k�;5�M�Tc����	r[�z{<9��K��'L�k�Ӯ�g0MeA|}b�[���9U��O%<���uF|m�tz�� (�G�g��)�N����{ź���#�ϲ��yup.�oֆ��F��,���4 #� ��_ �o���&a��,��y���9���Q	�d�w�Σ����U����9��6z���dBɊ�ڼs,�L@�i�(c�=��1jijӖ�x����j3�,7{���|�W��6�W��1��+%;��WD����3����5pgW�ZU&�2��Z�]i�
Fŭ��+"�v8V6�5�_��D�:]v��
�͋]��r�Q��W!?�wL��-VY��(4��#���ݫ�{U�6��z��V��!�:CVK�1����"5hG��P_&J�F,N| �?^��@0v����1�VPCV���3�dU5]ZZ65TC�Y�?�RT�s�9�FU�/�L�:�R��T�/L� ��4׍LB�8��V�eZ����'�6�E3_o|��L�W�5���Ԧ
̒�@7��N���B�����N�NEZv@����H'�"��U΃[���>�Q1�[I��y��v���/�Q���>�n܂�pL�%��M�x��.���E��f��,n�Y�R��Q?�?3�%6�(6���|}g�j�G-k&�n��\m!��p4a��Q�����} �yy� 1�s�����;jalen�xu����mLܟ��6��=7\A��q����6V�_���㻲���f|8f�q��ÞQ�=�c�<�ۮ�����tU	�e���M���
~|�m���wߑ��yh������U/�'C������B�CB%�KXlf�F%+شj���)�Fs�C���g�ESo�am�_�b�M89�~�u^����0#�=���gb��g����F�Ϯ�?X":���x��ǈ�q��jH{!�m�Mh$���С%?T��H ����ì{��Bڞ�A^C��2�e�j_����5����mJ���j)�kҐfeٞVk�ݢ"8��_��\�)�Y1�;>��uS.|��l��b��C��%�W$DI�hl���z�M(X��z�K���f@?!HbQJ-�O�}{����#e��I�#R-<���Y�i#���E�B�;�����Mp�4�A�k/Eau��ߣ|�)�2�?�� �!^r�Z��ȸ�!Q<s-�����G�k��43�j����逘�^{����e���� e� Z-,�| �䩣�C�.������sZ��~��^�����*00a@�p�;=�џ��t.����15v��{����;��0U�]b�Ĺ|pͰ�.Zē�I)���F�U=dÖzw�5��_	����?v�>;ێ?�l]�nǲ=�F���j�f��X}D}=�V��
 Z��6'�q��pN91��Y[�r�Xˀ��4aV�TzQ��7���h��QC񹘌ZO�	4�{z?�F6x�su��\��J��z�eA-���拚*&��@��9>n��"oD8oB�wLA���D���`�R&���u<}�׊�BH��(����p�,N�(;�#F_�T6�u �"��C�?W���uE��\4:�i��׼}�J6��a�y�����y��c��t_��@;�N
6��� ���m�c��ҟ�?&ї�����Ŗs^H�[#�8��=s�ޞ5^a��N�[js�,%
�ܿ�0�V� ���~[A��J��n�ZG�~S������Jb[�b�7M�S0��ht����-A��H7�(Qr�Ϭ�~Xx�&^�1������?2�dZ1�5l(��e@(���̧��G���9,��'L�=,L,�0C7�`t=6� ���A�ЛH�����4�;!��	����z���P��;��V.��
l�����!��_ıB�L�'�Y����A�����dL��.�v=�����ٹ�I$X�ٔ��p���:Vӷ_Q�vP-rĊk������>��*�?�/t��3G�ȗH�<��yO���+��/�т�m�(�������p�����;��Ji�fϣD_^c%(O�(�W�A���-ѱ�v�O�i7�Qz+�G��ڜ�g���jE�����W(Q2� ���.�u��e��(d�º��)0hks�0��|D�4?��{�x��,��� H�H&u����_��*�J���j5�}���i�c�OeJ�olZy=�Q�A=Uh9��s�g^�=G�t1��AQ
�O��*�CR��y�gߚbQL.)��|�m����\f�[S����mL�蠿�n�j�����?6V�͢���ѼU�Ê�>�>��l�k#�A�H*�qwF������BXH��j���<����i�G�������j�-�T,�,dr4��1=�����Z��H���ŴH~��潁�/�Z`/T3�BD�p\�L+s�ԥd���D��nk0A��v\?2&���)�n�x��ԅ:�T*�q#�YJO}3���/E��$^g��1�,��浇����I=NV��O���x�-����g�pO$��R�/�u>���P�ψ@��[)����a�9:5�$*7n��Y,.�#��@�LM�5������m������x(Ls��9���sh����j��8�X74}�e����A���N�
őUD		�98�R�5X}Lۨ�m'"@�6��ȱ��p1 m��"Ү&Z�tj��JJo�s}�? ���&�HmG�s�3f�C��o� e"���{а���\Cm#��n��IN�g��޾`�Za$G����]v�b�v�H���B,	r/NB8ֺ��*6�(W�r���h���G"��./�rB�a_8ed�*JȋH�WWe������Ǔ�z�e�a�.YܘMO!���U.C����YiH�Π]�r��^��*~�\��/�;�(�fߑ�`Z�$*�h!I�/0���ɉfq��#T�z��B�T�Au��HwF�##����+CK�`n<�"Ę�rlW����☃�!X�d����|߷����MiƑ�O�-���y��d@e`�.V��/0u��f16К�	U�����T�k�*]�`zt��{�h�t��������D��:e��F�j�2Eƌ#��T����
��>#CN��"#EE-�>G�cJY���3(��NR�M�k؛��j�����{��Ob� vA0��y��J�[�T����x"G#V�����9���Gv�P}o�,g3���S�fc��^��+�L�HG�F��.�����B����؂P�&���&���,�{�=c&���D��7F����y�rUW@)mGF��@�ɗz8:.��y��+\��"��.��D�r���Z��ȁ��2e�%-���{L�=��"%2��%@��ǔkM���jb��?���W�͕���5��m/·وc���#N���B��&��}���Gzf�2��HX�w��g�j���Ӱ�D ���9�"�?%�W����������B�O�t���~ <"��L%�l��fAֿ����T�{.W�R�Gn%^u���M3�6��p}��v�b�U��ķ���7��L7��u5lؓ��"	ʷ�����k
a�$��� C
�/7S�)#�T 5Q���3~��q!9�hDc%��>8n����"�J���3�u�YY�'�c��e�N��A�㱝���v	~*++�E>�M�[iY�_�2��YH�aD�D���S���akvUy㍜o��@)�CF�K�B2���.-?ʽ�|����¬��Š��M�����5 �.����;LgF坭K�E�F��ymu1���$�4���|h�����PE4D:�
@�����&��	3p�O7�U�U��C�K
�`6A1q/���EG�aZGwf���<�qr:��o��{�l�a �R7ٞKW��s�v�pN����n�,�������{�ej��#X=�NEQ5c����6189���_aZ`��V�e�F
�#�q����g.��!����.Bi	��3�]*�����#������ֻG�2�k�N�I��>��@2��i�.$��F����u5�;9M��$�n8�d�4�qRJ%��t(������8�`�D6���MN�a�:��t��^U���������4ˏK$�+�v~�b�~�Z�0�����:�Ң�����)*hΈt��
�ς9�EU`�2�<K���}��u�g&;�80��;�+1�OsMS\�5�rUE��?�K�a<��&�:4ƃ��kK���o�/���"��2YUL�cGCA���E�'z�l�Gִ��q��m�<��(3y煾����~�	VÐ�xqQ�IX�9ƞ��LQōZW��l7Mō�%��ׇ�^�ð�
��"��rqX��M81�����}�:��xR�ܽ5�Br���>�~���J�t����ea��sC~bU��!�ㆊYm�;�`�w�K�D���4r�K6��*r�[�&��F?,��Z�:����+��|��q�����G�hK�3=%������L!�z��������]Dy���b��J�s����m�3��H�3�%t�GW�.�����Ì�{�����6tl��.Pv�h��ҽXL'k���X�mo�=���z>�ܰzQ��M5�m!���v47 qn�X�w{�Q���Ԁ{�<�ǽ�22�TkX��	z�x�$a��x'��-��>P�;���s�˕aY�z+-�u���X6f˲+ á6翾}�r���5%R���/����#��B�������R�{$�jG#�\��^��:m㩞�T8��f�:X ��h����k��޶�[�&�,� 	ol�����@�dXv/>g�T����YxMϳ�e��=�L��\��_+�n���T�,�\�v�*��A��6}�Z�V��6����[��6SX��L��H��G\g�@o�=��Ce1��e��b�mb��c���E��Q�vUү!�j��i�[�T�r�p7lJ�{
@Xq����]W�H������yo����>Е�.�T���(���z%�^�O����p��p���Y�JI9�����9� ȀKXwB(V���0F�,�KM?���<7�}.�a��&EN�G��졘��8]�ԩ�*�)z��'gM��54�B�|B������D��2<�r�q�Tv�N�����g�E�S��������uWk���~�=���k/��-��P@��n�j�0�2���We(^�^�I�[[�NQ�9ؚ�Z�h�sȠ�����~m�Ȅ���@��?i F��uL��ig&Z��V��c�O=	05�ͮ'�{{9ne��ؿ�z��>y�H��B���Ԏ)�bﶀ�F�� JR��Y�R\qY����3(a;�&:Q��Jb_�{�Hї�9���
���<\�����8u:��Hf�Z�I��Y�3ʲ�l�{l��~OZ�M���{�a:�脀�|��%����Qdn�9��V�3�\�Ҭ��7i��A�XWt�8�P2!Y1�"+-G��"�e��w���јdC�p�*YDT��� K�N��	�w�b��EƮ�c���8�J���C4�ǀ�2�_�FZ���:܈���Н!�mֿ[dKV��pa��%�6G�`��Η@��q��͋�\�KT�y����X3=i��}#%��H�R�F�B5�Wh��K�-E)�����ٟ+��=_�7�o)`*�k�y��n�N�Ư")���"��)�U7��,��
��E�� Xud���>I�w#l-u,�O�pɌo��=Q*d$����N�5�L���&���2�$eN:�`-�_/�/|�f�X�J��%�?��Bs�D�1���x��D|�fw�c���IH��J���d�{5���J"2��( g8��E����=�D��κh3���{��"3�(23#�{��\�'���* #%nq <!�uc�K�qS}��FI�6<9��`���w&:�fQ$����0�;�V�RyIh�B!ݫάB��H��We	��E<w��\�<Z��X�M���u����:i(~|#�nu�<J���I��_��?�vYUڏ��S�]AiD��S�(p3�6��&
mZL�
a\j!���-7m4�jF�-��g2N�ż�:S *c\�� �C:�^�|�n$6�R����������pB��b���4{���X��]�X_�ԍ�PC��18������F��P�2���T�����|i�k',`).��ͱ���D}s���(8�'_R)�B��� !ԍ�����X`��كiA^5p��Ċ�\m<%�|jÊ(�f�@�ȍ*�����t��S8cJ��\�
!�x: ��PE���y���}�@�azd�G���͗n�Q�?�@˫Īsף\�(8�O�Ѽ	��g4�bK�z���`�r���4���$�foEȼ?���8�'|0M�%��,CM�0����K�L	����_Pc����s�~ԧT_ƶ��a���Fa2����K����d�MR�
�0I0�k��Q��I�7���p(v���N�(�K��Nȴu�03N��k�`�o I�q�&_���j�\̓�g"����݈��H]W����5��'J*�'b�Ҕ����Ժ��3���i����N^Y����A�"��E�	y�{��S�F@󏃗�.�n�`w`� V��ektaUy	>K�p�������X7*U�`��Ϥw	m4�A���r�(�2П˒$1�3�}����V9^�y��N�͈�V�
�t�A}6}U�)�K�M���0ucQ�m�N�^���N����0͝���h�va���.HU;n;�Μ����R��1�;4������w���&Θ�ޘ�џ@+�z�Uo-�b-�o��JQ��@���^���M��oG�2�v'�@�;)MR���,��.\V��/�>
������������"~3��":��_�� �Z%��2nK�ͭ5�/�4U�H1=9Nܭ=kÅF2�$�]	�Q�`�I���D�J*o!��{���ʥ=B �����P3]� l��J��C!Q�g�)|���N�G&��Px)��M��^�9\ȇT���_�3&5��0$��`��=w��E��~M�d��4�"��̡���G{�ȰR�1޹v����h24F����!}l|�oLo�6	bLV@`��b���ۥWGyN�Z��T��^4��}.�w(��F���F�Hsԁ?�[���\��J9,h�T�U���;},8Z��!����(D�ƅk��D�c�4N�ƥ��@S?v��W<ŉ+�#� �#'��?̚�MZ!�^m`�t�?Vk[�y���Z*�'g�#�����Kb^��Ǥк���0�Q#?�5 �"J�O@��e�XF�+1[��:�r���w�%<u�|��N=�^(�%]���)�����/\�C�T-�Zg�ϣ�Ӯ���r��@k�
�|H�]_6(�Ś"�t��9���+X�bW����������������/��Ah�}��!�T�~� _a��{��ŀ�.��c�d�@?��%7����t�L��������v����l_�����ٞ@��-���\�)
(ڊ?�OswĲn6�V|d^i��7��α�D�UՐ��,�m���<� �my���py�N�
�^1���&@U[�y�qm\Q�`��Cj+��W���ty�uI�ye�c��0sk�׸�+�SaX0����t�z��by�X
�F=��F������E��F�:��v�j���(	��  ���vn���j|
�ύ��\Ň�"��@��b �z�0j���ER���º��`�%�1�tjI8�������P6{�E��L`Nq���O��o�SѮMOL�\4�lS,-H;�|I/ø�*������UwK�6z^��Ŀ�&���z>������1 ]�~���3Gy$�:s�s��5n� � ?�+w��h$`����.
Mb��X�g@��K�3����ҳ?Soj?j&<,�6��T1�F�	�,z%�@H*Y �����t �$��!W�}��u�� ����J>{�ފF _�1'���6%T��8bZ�zKHv0.�`Pz|�WN��W��D�qʣ�w�ʃ����+��'Ms�����+!
5x�ü��VG/�Z�*�(;�e?�m{��s�h��=p;��2��u⠾�x�fU#����⳧,��K�~��9}[:� ���CA+�%/�
e���n�)�*68T���?�I_�-T=�W��<'���X���A��6��9�s�皈c�H��~,"��vj��n����8DP~o9���̠��&��+g�Tګ��*&e.���H>c�o��0�;�O�3k���-և�/�4@O��+���Y��J�DX�zv}'��<��
W]�6��yF	����z��[��2�dA��lab���FzW�ۣC����<m~8i.zqj�	�Hn�>�O�H�*"����U��ّ0��\��b|C��$Q��+�K'Z�@���H0@D�I-cp�1�3�1�O���
w��<gU�����#�J6�W����E�#Ҩ��T1xF��>�JC�v���5]��a,��/�{o���h)y�nD��xE;�}�[N�h����PÄ�L&i�3wZ��@�Ap��$4����(��M�}1�I~ �{&"v^hL䞳�~D��5�E�nu���� F�c���Js��P^VtFܣўI�ư);r[���Qn	A���� 㭷��0jE?���H�3��z8[�A�#�����-}�R���4�0�.DW��ץ^���Dv5���;�5��YT2����mw/G���N�c姷d3���̈�m�5.w���i�}F��c��{���<'24�r.�=�n%�:W(m��-�Z����Ϋ��Ί�&�X�Q�Ua�C�-�c-�Գ��%�O]�� ���2��Ӣ�������%�r����_rW%���^e�N�Xbr1���"u<��h2��*S`A�q՞+F,�]	.���w�u��Z�epz������^��$�Br+�-_%�Kz�:V��w�J�^R�n.҅.A�w�m�������Z�����GiI�:����q�g��������gX30� �/�2j�Y�2gmPj���(M�&������Jo;�J�Fr��!{��`o򸗜�X��{�Bd����?�H�%��n�,�;�.�MM��@����iY�3��ʙ��}OpH�8�y$�0�Z5��c�W�z<�šE���/�,�96�W~��o0vg�2����"����k�G}��3����������19F�%��}�1���Ƙp1_/�|VrϤH�O��QBb���d�p�^9�`;�S��x�5�0��]��7�8��rD�pn-�Vd�N������9Ϯ���X_�
���?��V^%:�:d�@�6.�w��O��V�3<Zb>�`��W����G�Z��m2���ȬcA�Yg�������%"h��?D�bm�����[�I4f�4_~��:�!#�~���o�JH��nS����4�ބ�� _�aI`��:��;z�7��#m5�J\D��Cc��J���S[�vEb�4��$ ¸��ܪ� ��[c�Y�J���[eد�B�
���|�-�-�Y�1w��<��J�Ѳ�=8�#�Y�G�����&�H����2��)p����i����rNm�Su�D�<qW��	:O*: ۬kx��|�l���n��0){|����m�餲��v��8��!�JH둭�` ��_�O[۠�ޔ��_侂l!����C��Dg�q�{��� ��?��kȂPJzQ~7�a��Ě��/��l%��*N06V�&��y�(7���1�z�y�:8�Bh�H�0�	��^��X�!�\�n���J���/��KWV�a��KϴV1.�:K{I�2���Nj	�:�����f����]�wS��6�?�D�P��=n[:pҡw�z��6F:q�����+=��Y�k�9���m�E�6��)��(x��;߶H)Š���3�`V%8$tcy3�8;
�yL֥Qf� �j��8T��}�qc������,�R!�e�R�mB�OT
#�8������]�����~wx�	�R���^���*G B%P�Vz���O�EY���6~�����vgC��kCp�`xh�ݞ�vВ�_�B�!�C��Q)l���'vvӪFU��jgqT�[9�0z���b=aH-V`�zŗ�H�TP�bGND�wڕ���ۈv�#���A�TXKX�i,qM�))#J�m@x�r��v��p��U��bYt��B�P��s������Ǖ�f�U�ڋ�GF���+%������*Vb}�K}]xӆ"f�~,	����e��F���L��E;�w�x�N�����	���q��ij骔�[i���Ó�]Np��:�Q���ߐ���k�*9�Ly�#����z
��]Y��K+���	�ӽ �C���t������w8#�X6��߅��B���(�t�{�yqqթ#���9�k���ؘ�3r�́Z�nx���1k����������i9�<�"/��,��p�#U����V1�ߛ�<!�k6 �C�Ut���;=Y����g��n�P~�g�K�i��k�{2��S��׻&�))�U������� � �(�zKˡ���+ǲ�㩡�qCJ�Ù�>� �3/Q�Jo9�u8�ꀪ5@#�a�a���xQyp����@08�oLI��M�����G��##��D?�Ψ�4mZ+V�u��]���h�^))�1E�4�"�~C}��Ԡ�h(�>$l\�/�ɗ���U�?�!�4�lV+���%����}�p/Sq�l
,�,�#ܜL����tO��:�������l��H��� ������R��䐤�{/;f���*��>�9o��u�c�j�M��/�
t{���C�B�Ό�D�_\NR$���$F~��*zY�'B�
%�<��%��;����y�5� ����Sdeh
�*�$�-���t&�ǥ�ZT]�����t��qi��_��E�#�8fC`G��N��jy�:�47�p�X�6��DN������i��"ߒ��X1�*n�Ts�+�G����9IǗ�wA�wq�����ٲD���驴]��?�>�ȝ���YL�b�;��JJ�A�kW�Y՜쉸�-n�**b��e�m���;Lm܌�M��[w����XHlw��ߪ=���%C�ۚL���������Y*O��fѼ}�/
�ϓ�Ds��6�qD\�A��0
�L�-���`��|h��o�:)�O~P��9"���\�{N�U�{ѐ��f�p�v^��S�C��}��i�X���(FQq4%�%�X6��i��y�>A��m���}�9��ڼx�l�};�VC0�"'_ܩ��rypYN!W:V��d|�$�c;�Z輓�<���/d�(� �̼�8���y�Ob6b?�n]����X*F�O���p
�O��V8��=0�����о|�\����o&�a�0��l�}D���9�T1'�I�����>0��Qzэ�){�� �FJ@�j�[����,��n�]F������{�uJU<ڴv5�w�&�U}Į������2�����(���N�νNB�L�����aq�*R\����(3[A��4�$��E��x*�q�h���j��1s4<��i�^��
�a7ƺv�D'D7i�,7���
�g˳�{ҩ�e.����8�?��9��R?�!�6}ݹR׹:�5�(W��7`i�9w���>��^�Y�T,Kyv�o�=�+�,C�4 Zѡ�DP� \�		������A6��^���i d�qQ�)�3���1�&��U�HWI?dj?Nq�>�\m�y��)>Oq�G��{)�<�J0��y��*��:(�Ft�A�������~G����i9�[�	��6����m9Q���	4=qr4Z�\w&?HUd>��(TWX���&l��Ԓ��u�K>��| �I��^P�j������ȧQ���9��=l��H1��ڴjY%W����o�0l�XR{/V�7��}��ޕn�h|�xU�ރ ޸|c����'�'�λ�o�d⵲��;��sf=ܼC�G�!�àls���N_?-�l9�U��3�$D|*���'"ZR��*F�Ӏ��=o.�Ŏ�Y�I�*��G�!ڡ���$�ր���s��/zN7FSK31�7���s'�\ӌY�u���;�u2�&L�>4�4��@�M|L���1������P0� ����6����W~�n��E*qL+Tݚ�~6�&дF��t�淪����{H����Nl�"b|�ڻ���Rh�:j�G���m�]h�c�#_s�<z_�����a��.��T�w(<�C^�j8C��>�2�mG���a���� {��^x��]휙���^�	�PmG���:�ᯫ��y�I���P	���s'�Z̙�~F֟1(:�݀���U3x����r.##�;ן�;��*G�q<\ߜ��M��+lws��3�(33#��0��W\?ƧA�����i�VF�����˘t�J^�sFJ(��#O�u��+��&XA8��?���G�p��SI��כX�Hb�!W5��7m.��^8�&�6�Rg�d�t&1a��;��I�r
���L�P�(����Ϛ���.Ⱏ}�^c`j�(+l�]<�`�F���<���4�w�=�y�j3�ጺ�5i�է9LG�����Q��qxF:�x�l3�@�����������b��%���Fm�b�;�#����Z�D����Lo�2�2t�Y�*��|;~c���lA~w�m�~+�1&	ɯ��4�BJ���	I��{����}�j_������7���Mer�~�5 �&��ݺ�9v�_݂�FYj=	p� �DA�~w'��#l�ȱ�xJ��Ϥ�l���Փf���V�@�7c��FO%�O�	�R$bk��
�-йM�o��� \�$3Pa�h�Ev�m�!�,d�"f���-���!Ne��-���{��H[���G����!1��x��4g�����I��j�j|V�$�V��6/e�jC�VN	�9e��q]I�L�kR\���~�:n��	ldӄ�{�8���灊���}*2i^��W�im���y��T�=c�1�=n�[ĭ[�3��T�,��7�i�n��Z�:dgg��ʴ�0���7t��_~>b.�վ�)�u=.�Pq�"��r�"�x�ʛ9�P7Ȃ���+��q�p�)vesH\�
��(�%�����Tz����ѩ���2�*Hkk��W2�}�9Rb�w���x�p]oa���w61�����#�~2c?-���Y	�"2��Y��:K�u���"!�7�r�6?V�+�������"���a+�Y�T	��&����.:	ES�j��:;��^��ϝ�^9�(�1h�e��j����؅�Aj��mnyLYaDֽ����5�*���6���ڝ�2��b~�m�P�^���x��O�Өc�84%�@��
xZ�k�B�7n��%�/�����} ;ҋNɬ��^����Ϯ�h�"�쵩x�k;ʵԷ����P�vc�l*�D*i=�Ĵ�,�_��?q��ʜ�(������RB�ް,0��$YY
<B�X��	C���f��m�R�a�C���D����Y�*�{��A@�C�p���l8�˜�+���q���H��/��@Xm'0��*����2hJ�$>�5$ja��R��y�w2��~n��x'�/WwLf>��W�o���>�&�o�)�Q��:��:)�[�����Z�t ���a�؇Q]�.��B��h�ّa<Oq�΃(����O�%N�MU��[A�ʠA���gJ��v�b릜��v�;��lL�I��{�n	G��ˁ��H�G���{n�s늹��F�J����K�VTED|ݦ���8�|�1��	�T1�YLc���O������q5��a�#��/EW��\6к�lA���f;}��M���K��c$�V�|�5M��G8{����&5��ɢSgk/�1�����j$d�ٮz���1���=�i�a������ �������1�j�WĲ�M�������𻋷b^tE�T)ـ�����Р\�~���)�X��z켳�G��`���}5�Y���//��M�Q�B�6Q�z���n���'�����t���Mk�l��n{�lf�<Aplz3���e��O��l3�B�:5�TI�)N�"|ΥEls�O�	���#`�֊T���������_�Eׁ���C�6�5���<^�����ֿщ	�6i�u!Y���>N����J��+��q�Ĕ���d��}�u#�mhy�W�࢖��Rm�9^2;I~gcK��
���2�����R�u�+�C,ށn���",��=d�X�&������XE��d�tM`����~�4):������>��+��i�v���k(v���A5~��;���Se%��Bq@�U?fLγ{��o)�7�9��y%ٓ)R��j��=�m#�&�5��6y1�0�N��f�o:gdOщP�3��K�޾�z%�M�o��h�
�7n�u
s�0
�����`0rh�&���t��Q�� ��F��Zc���|]b�U;Ç_�,���+�ɔY�9+���n�{��^�$���V�[���~��M�熌��_6���LA������hi�a����{@5����Y�GA�L�쿼�]�����6�7�=wN�E�|�/:���2SY�$eZK���i�fl��hkCD���Z�����_M%�UZG��8���sr����T�ʫϗ�i��pZ:�z�Ƀ�����Q�E�.�0��<� g�P�F��1���!���8
�B�ӶJ?�T��l:9G^F���J�1�#���#mM�|����o���z�k)�uIo�F�iɕd7y������QHBx;��Qj��~��K~�0KD�s�ҝa�g�޳�E~�(�����XۚÔ�?��c��[Nz�v�K����^~��#���v���^� �Ǯ�ן�����:�*6ǣO2�8＞Jy�/� ���}��z�{�bl4���"���y}]G�.d����i�w��i^����@�gYͦ�b�~��gt���莯��@�?T6{�`�uH ůE�̺��6��H
q	@۔��Ǟ���aY#(\Q���D��>}�&�pi&_1����ª�nv����N
[��0K����e�\#�u+3�{�1�}yPo;�b�Ҿ���#���7����rf`�#Il*���|��8�]G�𐥞+�)�Ϻ�l��8���$�<#빳��)ރ�k�&��0�H݃ˑu�#��{�8�nd=t�@���#?v�p�w�i	;� �#��g�o�DẔ�E"lP<�L���5?:	��k�A*ȓ�e}$���#a7���ct|�D����I�(�T?F�y%�OxU5ŰEC�(ztO��X��gg
vV��H畠�@�;Y�m%����j@�褺��`8}v,L�5�XUN[����;�8���F�^%�̹�D�l��0�<8OL�d78�7j��k������=bƲ�cs+�iӈ�l+�|rf�1�U?����sUF�7�&�B�W��Ip��d��P�mv���b���oX�_���U�yn����r��P~e����I�f�_�"����p�Dp�z�o�\h���mFX���������T�vV�3���u?Q@�L��H
�k
}~�^��2��m��6�F�.��e�"�MH�����3��*�=�@��F�r�I��a/���� �䏔��7�MF�ˍ_����^�p�O�J�e�v�U^[;y�\�K��Gc����nH>�fĿ~�A��<�5�]��Rr"<ȇjr�/��'��@T�T�|�z�w���j���_��Arc�'�38UE2��4`=����g[q^k3�=�%�m��݂Q�qQm~5'So�"f�x'�nyb�s�����S]G�\UΗ\��*�,f�T~]d��H�h���/@I!�5n1p��9���8�z��m�B!w�P�5� Oe�$��.�W"n��@;s��ר%�e��,*5:����vJ�#vH3`Fx�-�#wu�ѝ4d=���O�=M0�;�O��CZ���|��q5�*�B(�W��V�wz*�'Tr�y�{��cm��N���%�Q��Zy�v��@�T��-Q|�6����C?hF�JQ*
B�5w�C2�55*A{�vq����~��l|X�?,�Mvn��)��]�I?H�|�2��E,ڛ�u3=o���8Mb9vФ͞1��05����� �� w+�f�^����ƦM�h��m0�;�C@�=8���%V}�R�<�ׂR�G����� ͌�IK�L�����\��9a���s5:��[t��Ȋ��*���}qNWƄ�jW����9�=]�Q�;z��{B
Ȗl��܁ ���t�5x��C�A=�-"�L9kt'x"	#�Fj�ա�i����z�9�
@V�?!��/�_��u�"��*E�m�N>�s?��)��ڔ�:t>����3oeS�a��5 ��@������i�J�z$�R�x݃��V�i� Fv��  �����YN�����^�����sh�!���+�*I2>���CeO ��AU F{���]f����9@����s&zH ׮1nn��A~ʁ�L��݅S��W7H�����ӈ���f$�x�M��t��pL�T��L�RH\P&��#��@lv��I[uu�	��Uݾ�M���n�-)TE��t),�sk~
���m�ݑ��������y�5�#Ԋ�a�*oQQ�v�Yiy\�
OlbR���wEH�U'Ԯ{�`�\�O�pO�y��"/FСe�D���H���$��bR�b�"�����o�#MĎ��@�(⺪^���a�w@P5�'N0���Y!��Ƒ=�ٷ�Tw����:��:6D�&�kZx,!��vi�����4�[_Vq��7as���e��$�^�]�q��'�q�� �T�\EH���� ��Kb�J��q����[�R��B�R�[�2�3eF������/����>IS�"��Y�aDF��S�i]ځf�Ys��B�.����7��9��/�H���#��y��7Wm��'��X�o��t�0�dȐ�Z���,f�������G�>[u���Am=�-W��IpOK����y�
�B�hJ� �w��h�&,��o9�$
��T�坌%�c�;3�y����WOĜ�������:"xZi)?�չ������XԎ �`*��~����wk��J�]��-�P� ��9u(�3�5�B������ �%V�/��ۘ5R�o�b�N)8�@���[UA$��.,�';��<Xl�<�ZJ46SB��gr��cLI3�C�h����+�gn����������o����I����\����l# �4�������aʀ��Kj,��Z&溴�U�!r�LA,?�������5�YR:��$%����j��_�X��q�И�_��<�&@�����kp�3w��ي�>3|0������F�;�3�P��C���v�N��Ȏ�'�+ETƾ.h�*B����g�~H�	R��+��8����؜��q�m@a�P�m��t6��-^3 M-Z�5�ȧ��Dx�����J~�30g<9u;�\ݷ�ݧbu��a�3��2f������c��EPx}��I7]g�\u�6��X����OHP��SZ��ӃwӺ#���\�Za=a+N�
Jv���NVA ��łu�$t�����$t0*m*#���l*zHYz<<+��?�q`�&�
O�y�	:�b�s���
/�d��U�+
:m�c���ݐh�jhLW���|H�v���r���]�����QN5�22�}��#�������H�%ֿ��.%b֐�0 �����Zh�,s�!ɹ��Y}�3ė1KX���c�M����@����سFڠ��#�Z�� ���DR�Ù�Tz�f9�+9j9%�HVK,r ����L�)&[�MB��q�	(���&;��:��P����p�pwn�Q����-?k<����r�@�DU�srkG�[b�����76~����MMJ�ˉ�'Dq<,����$-ި����LkKP��OE/�<2�nW����0���v*H�<�6p�3Tp��+g�2�W���ͨ��|�y�Ȃ��G�O$�(|������y[5.�7�N.OƆ��+#h�3��\K��@��Q�ޭ�lȒ�����hMԬ'�ʰ�$A���o<j������g��ΰ"3W�FN���N+CS&��	/}*�L\�Yn,���"�o�P�6ze�}ծɣ����T�Ϭ��b����}�A�LH��kɁ��B�^fO�ěH�������g���>�^몵�FG�	�
�Q�|�W��|���u+��c��~�D�j1]/C/oj���	݉��v ��j{� �=�x$�����Ĭ�w�4�r�����G�a�:L�O�A}�Jh(~�h��S�d�>>I�=,��	l.�Y3�9xC��>ք�����?&�~������rp�9���t*�6�ڨ� B�Z��!�-�7� e����oCq-�#���7��0�9�C��^V�
��.�v"8�P藐������GtK_8QJ�L��*^�5^�T3��ş���A���Sˍ�fB7�ݙ�e�m���@S�bp�l>��Z������h�,0���b(XI��j�fuɗC�d�J��E/O�nc<����v�
���m�I�z:����C3c^������1�g����oEQKS �<չ�ֆ7�$0i��HVH�m���<�pF� VِNw��v8%�{W&�}e7q��p"۪��~��E����k�
�m5q]_]�F��,C���)uM6�3	��b���t�T��A��bR�7:r+w�T-Ȅ�0u@4���\zN����0p�l�	�Z<T�?kl8y��i�6/�ܠ!P�<r �VK���Uu�'�����T8#�DP�c9~�m���?2뚣@pa�І�ln���+XwG����f���N���+�!SJd�L�v��;�]�`��Ȕ����ǳk�rj4�k(�fF�M<��K�O�O�O<�M�
�|q+z�L�3��t�a�mxД�������1F��?��QsI���B����#�_���X�8���[���:4��qX�v�Y��Oʙ�W�q]R`N��g�q�a�^5��8�/�Kl�; �T��-v&%ȱ8��A�p�ǀ�r��G��Q�U|�'�čv�諘1�� �����!�:��Z,6��}:��j�>�.�k��ďбB�p�x�l2���C�©T���l[�܅/m�9����љ	�1!q�T�.|���O;����_�^[���h�; )]�U(�OŴ+��Vm�W7���| |5.���\>�q�sLfD�;M;uM�g4O=�
?[!�W�a�F+�}0�G�1Vm4{��x,O�U�2�6����������|q�&�� �d�ڡ��J��WJ�3�����?���0X�a�fr�߂V)�.ɢY�1b{B�$Q9QEȷ��M���G3hl�DY ��;KtcӖ��͢`�wggkU��'\���嚺��珐S���7�3*ە;)E���<<��d�܇S��͚����9:�t������p��QAh�1~g�J*������ ���� 7c�d`�ן���GO���yw�:�b�WyF��7B��}*�P�{�ho}�^J��W��X�Ӵ�S5 @V���Y�$�hv��BJ>sk����@cu�!J�#-��^c��TNn�w��ȏ�H��c�H�_��o�=��oq�����!��R��!����NT�|A���^���4uIմ��v��B�m䗱��f�<���+�	�"�FPTe��px<:��巤$���FJ7�����$�#��.��̠}��^+�8P���2��a����p4Úp%�g����obOc�	�ƫ�Q���N�P��aأx6��hE��O������.���*�1�k:qw*dߤ7J�(B���m���Q|f�gk���{�4��YݪP�W��9$���_Yu���;�P�^][l)j33�
:(��9���J�3�͡O�Rj'&��D��jηl��Õ0gf?1��ʢ@p�J�m��D�H��<�|4 �(<���Hh��]]���Ϸ!�J(�o�"F�wIC�Μ����N�75����U��ӷ�y�xğ������%�"cs_'E���x��[R��І�R�3�v�4�3֛[<�l�u2�6){�}{�zu#L�M��p��	"�� �)9�����6=�4���;`��P��DO��x�l^T#� ]��e����s}^]�A�^�e��$0�p�L!~���_A#����+�*�p�����a��Ag�Q4 q�C�0��;a1ݖ�2�@�GL�NU�cd�TFki��"�i���!�!a�4�~����'7us��e�Y*
U?�J���.�|��0�8h���l.��~����Ӫ���@����QT�/��L:�b:�d|-K�,���-���Bۘ*��Q�"�M��;x���,̔NC�4u���Jp�j���i%�oi��ͪj���"C��%�s��Zf�a�W[�b#+��L���?���Z�)
�_���B(�ݠ�6�@��M�=�@N��	#ۧ�)��ؾ9��^[�T��q��|����_�õ�lA�i�	|{�}��*%}/4jRP8pQ��S���Q���l��'m��Kc#��e5+�Y?F@@���wgeG��L�hh�+*�o�7 �kx�n��o�R2Z�T4�f��"v�Y��B�q �@`��l;U|dݖ
� _tE�Y�R͆cKF=6ż��-ʿƗ���W��/.
��Q�Vy	,"i��w��z���� ֳ�`?�8i�T���)�T\!�Hy�=��3��Nó��m�w���ێ�Fu;��J�o��u3@��[�t�����˰��P���gѢ�K�;ʮ�<e�5T$�M���¡�W��A��2Z��8!���j&;!��\?�̵�c��:J#��{g;�u:�E�#���I�%D�YŅGb�n5���D������ʭ�H�t��� �f�6_�������Fr(�����F���7?V?Z%!sM��I��Z�|�up
gr���un���A�d��搀�[��TƉ�0$�����ĊQF��nR4G���C�[��g�킮����x��E�0��Pփa=��?�k&inf�k\�*WnZ$�yhg� �k%��.�ʖz�I�44���u���a�5#���Gy�,G�L��+�v}pl-ys��$-h�=E¶"�l�$����d�e9�i=UèL���	����4���*֫�v璠�;�Hp�n
�Ol���'n�YxTWUS�#V��A��)_�
�<�W��w)��d�7F��g���
��9��°>�Y�L81��z!=k}���J��6��8Z���*����Y��n?dU�˥��	:���P&���C����mu�^m"C.`�4��Mp����5���U�
i�t�o�8N�Rf���4�0Q�VyX��R������s�V紓Lw��Z`��Tt�)�٦�}�qsFVE}~��Q|@�h�aW��:�����[a�Y{D��������*�q+ЎO<)��FM���9U{e
*��Zx:s�p2���H�/������bJ��F@A��&
&-0��{�nQ�Yю��`��cG�MU�s�dV���9���JF?����9kX����@���3-/��r�G�@>��Ih�m���u��?��g��X�A���=����@H.)�3��o��+Ԩ�̿�+4�M��v��X"y�N�6w�b"Z�4��pm�/��0���#'n��'O*'g�Ԏ.G��n�!�e�B|h6��?Q�0�<�z�Ȝa%�ɵ�Zj&_C�6�<�%ϊ��۱A�M̐�
F���c�u�~<�(̮������OJ�bf�>�V�@� �n�H$����x�te�#~�5qM1E��&�R̍�l��u`|C���t��z�1�O⭂{Q�6w�ԇ�;-Q�"M�=w\�ڄ߮x֑	-d��E���r\���+zk��=BZ	��M��x̝_�np�%#_�h�
)�^�8vB��E�͸�xߢ��
��U�~U��V�J�'@��Ӑ�����O8 չΑ��W�ﭜ���PQG��@���� %9���Ok���g��M����L��=6��u��@T�q�>z��@��?=@�]p�ck�˩���KK�L	��\C ����=5e�b��<��� V�NO�X�1AF	<�d9I�X'x�k��?*��+���e���kk7ڎ`*�����&�$[����s4�H9���GU����r�H� �N%oIy�e��0��������yfBn��Z'�Q~�-KμOC�����LB�	n ��FϸY�����q����\PCI��/X	tK�h���w��i�m���h��8�ŨE��`�R�3U��,UP(�ϳ $E�%ռ�N��O�SU�݇��+���z@G���pu2I}M�(�pn��7���$(�lɰ������Bm��㣺�דi�����A��]Nw�M�<vR�-L9��@g�x���T|חCb^�$���~*�~�1�@�z���JQ濦���A���6Jķ-�� ���tSy�|��Ь�ͣ�f(ꥨ}�s�<]�'�na�6p��<�6�Φ{cx'hJV�E<�7�B}?��G��qf���&()�Ű撝�U����H����$>d��h���3q��29��r�!�
M���K��������#	�1�x�?�������4QG�?�vQ�M�C���(�C������:h���s�b�5?��v"�UW�����}�"��&��ٻae��;%]��-���uw����ذ+++w^OQ�6�T���WӚ�������'1��
�������#���8����ai�֗O��f�ȼ-z���=M�׬�Ǣ�iG��Q�hPZ�֣T�e�`5����Ƃ%�AC+�GH'��V�ԓUD��;�B�����Q�!�ɋ����ѐڒЂ����Y��|22,�J���p�\v(��&E�9uIvU�yqr��`��4C�m��K,�m�4o�a������ �\�|T�&3���>̖
g:	�_{�����H�����&�Ĕ��N���[i����w���;�I{{>��%S��0 �3l뼕�D���"�IL�I�q�a�c�;�p�R0��'��ي��OK�)vv��:��.���R��ܱb�kv�l�	E#;�*nl��u3�����ģ�#���ɬ61�Ӻ1�(RS���Z�F��R�V0L}~��Ӓ��ZZ�ew��Swor��+i��V�]����U�ij���9� ��v�sZ���e8���+c�x#�%y�"٦4��Oj�"��cb��<o������ٶo�O��g�6.�a�m4�s?nAҧ(�������b;RRT�`u�1؄�0��'�+
��Ot�q�d�R)�$�yN��4��)@�Ը#: Cq!Z/	�^�yS���T���ŭq��UP�J�Gy"�ޡ7�&���&L��+șj����Q0�pލj���Y�؝�6��f�;��l����)u��pZ1�?��c,f�d2�f�:����B<��ì�]	�ێ5NG�����&�Ed',M0�N��s��F��.d$lz0�u�Ǟ�����W�z��(C�[�	�����?l{���|�szҙ&������!	0s�{��PB���GAB�ŭ~A��9BJ)un�"����B�<|K�?� ��䒲���P^<��Yt��2���D5�"���;'���=y�v���*��l�[ ~Ї(�wt>���恌3��N�'�m���p��\�h�2sc��� �H1�)�QE�؁�M�!N!G���=2ѱC�¸�^5�'ap�S3eI7coY���*��b�Ι�y`�ǯFg��Rm;��jڪb)�6���x����Pp��B�m�b[aY7��A��~p]�D ��Z���|�~�^����l�~9>j���$�g�Y�.��	����A�͍���|W7����Pc�����7�]7�`�>ޡ�[��gL����Q�l&��T��R̓~Q�f����u`��:�p����w���1+~�P.�S�VHdf[���.B��4�#�����;�EU�4䋲��|
���2�T���}_�7S�����t���X�U9�ana��.H��*؛]���Z/�!��ny�=��Nu�=�u���K��shcß,5�.[�_W��M�Z�j kZ�BY|봃@�[O��@K�Su�7v�Aw��A�տ6�в!�n�	�StJ
�9�v<����ӕ�a��#�/��qς�hO�*9��t�xmJc+t��	?�'�K�%y�V�扊	��2�N�0��rH*�e���1�ш� 8,�v!q�����H49 ��5+����O�Ɛ�1)`r��D3�17@yn������DW"Gaq�=#v�#��0Ɣ��r���ɸ��bOt��nt/"�]ae��y3bg�����Ҍ�����Z��'�-��k�*(n������]?J�Rp��Si=�ɠ7���I ���B�k�eM֎r^�ԇ75p�ӸO���+�;�g�^���b<v��WŁ���˭�W�s��\���� ۣ>�&�l��ڹ%	�mYF}a�J��Q���l^����
.�ֳ_�e^�n̳�S��9�ݰ������2���"�"�c��{�T�x�9�sZxE�����o2e�l����qXo�/���������wr����v����ue��"�!Gq%�j�db�c����iE�p�q0���7�U�VY ����k"�Lm+ʫ��Ԙ�������t�V���"�)bw��_K�8'����~��"	�=Gѽ�,=��T�}���P?���z�N�B���@�3��4>��G�.������&KB*�^�136]�M�2&oQ}8�&�AL�R���mƆ��\$�ǲf5�,O\4\x�G>�����L�i�,.���v���e�@�ܹ�z�UX��Ī��;�MM�`U�2@�n���z����Z>0#P?��)o:ʔfy;PG�,�	�=�=s�9ܢe�G�zę�c9�=)�.���r�H���`������{��r(�&���K����Q�;�$�N�db~]Z�b3 xW��(I�K1�PB�L��h�&�t�0hJ��u�g�v"�A>��$�{�!f���\:�7+>v6ߢ8F>'�U�
�%�S�.�H�S��^�֗M�Â�L�NX���6�:٘#�2��k��U���%���z��Y�س=�����'{H�^�`uۇK������U��h"�� F��(�>�v�3Y9ޠ+]�N|���c<��ѕ�ELz{x����� ���T��z�	�Z�xB޼S�.�� ��[Tm�Iڥ��%v�*i6�H���յ���b�k�|.��4
��6�ɛ���3���GE������L����&.ib����5k��7I�Q�[H����z�������e�}k�פ�y0֓���G9��� �L�L؉cc��t�Y��X�z/��W'o��h������7���6-��B�{����4s`���/��L�gP1�[gr��ݸ���i��ԞF㘏a�4�C�Ҳr#�r�(���)>�K��C��R�����&�j�C�)d���;|I����?�řa��v��n����,bY��գm��n��,�G�����h��-S?B���t�!�<owV@U��1��^�2�qk�}6���Ed�����b^F3�S�+�3Lu,P_�q�u�8=Jܻ�O�6)������)e�X�S%f>Z��y�����`}���x���Q)���au��xu@�����[�\�܌��U�p�|�?X�5H͡WW��䰠�h�C�b�N�_S�{�#���k𬉽�7��P�ޙ��Z��ِ�1e0O�nB�)�Ǌ�iᱥe���V��?MHS�]�ݤ��]ƥ��~� �m*�ʡ����/Y��O���&|XJ8fV����q����������%n�� ���%��ݴ���؇],�+�:2>ي�o	���0��OQ{0�E��)���� �<�^���^JW_7>/���ah�J� 9��>��k#�@�_��.<���Ҹ�+�����!WjRSC�W��0i|��q������R���"� 3h��CC]U�����9����E����p�������[C��e�Z����J�[2�D_|�fRb������{%�$�䚍EB�a�N�<��ᠩ�]%�~.T�x���[-Y��Jr�jI�>�'ݜ��s-4^7w�_��x�b�v+k�O��C���}96`6���k�W��Ɉ�ܷ�4�}���pq�f�7�b�9���|
Q8�Ғag�|ًl���Q�6��X��������|z�;n�ӱi���&�cG0�2�Sۢ�h9�wh���5~���]��;JIs�R�Z����:5������h�
ް[�K(�7:I�S�#>�ņ����A���{Jt�|�C>U�H<*u �����eX9��H��-�R��e�����[$��^��:��'�ZpIDX�g�2R�ޜ|����p��V���ח��倫�)�X����$7<��q3e�ـ\���+��I��	i�* �5�:��A��A��[�5�`��8ם9
?�	��QM%��I�ɾ(p��E���@��Ap�}ӷ�owgDM�����c�QM89�J��j'�lo�к\�j0ɪ]C����1�����9)(��C�H���&Q��f�5f�/V�'����C�����C�xb��p���(� �-
�i�-D[ِ���7��_�����:�?�`pQ�{@��8@�������F����_��=��|ٝ�ƻp �@��j�TDCao�B�?�#&=U���L�M	���B�4;�3!����R,:�Ko��M�B��V)���S+Y���C�����kvˠ���g�h?�R���;?#��9Εg��L~R]���d5$1n��9�����ZW|����V��]�y���YG!�k�m��`��&�*#~�E���G+Z8�F��C0	(P�������t�0�I)�s�A�W�+2�����C� F��[��}�~�Ց< >��kD�oY�z��cW��ҵ����J
�y�S�׀���ET�==*�O�
��m_�_S�4ΡD��ʹp^���I۸̶����D�֕y�f�:���$���mC��d�e��(� �v��dY�n����j1K�Y�[q��/b�C�x��)׻wqX|Мvx�.4m�����\[���Y��YE��}�A���3#���E�:"j(�_�� ���	�J�%3�$8��+��.����ۣ�~�om�48��{08�f��*3��
���=#�4��*��9�"�۰�/G�b����E�>+Z�ro�#k��'ӱd3^�9T�C�L��.`���a�A�
/v]�S��p�*8փ�C�<�y?1<p�*Ɣ~ǘ@������y��ױ�8���(�V����,ꉱ_Y/�`�"�Vxz\2"dyHsDC>n[;�n�*#�����̈��l��v�����辝���Yo�X�}!D����ol�y��4��='.��gƞ��Ұ��OȠ�	�#6t]zq�:�9�RY�a�W�$�}�b\o�}�0�,g ��R�݁0�@ t�o� ��DV31�����M"�s�l�K���	�'I^�g�Fr�iJ���K$�b�R�kvo�k1��t%�z"C]6��ƍh��
��W����‮@i����*H��vk����=�xb^VM�7M�2I�z�������o�UJ���҅��e�X�J4�"=z�qPۻ�Q02��X����
�?}8��~�[�浚��R���[�~nC�����2���VP�'�˲��h��[���`8��+C
�0+6"���B��%���&:t�^|�w��6!Y�7�'�Q�4H1�25:���k`o>�">\����¶�H�:#��|������њ�TC��{#�p7�M��]�����҄}w���$�#v�}E�+ݣ�2'f�}V��%Κ��lC�)��iQ���"�-<����wA"H6��-i�V�J��1S�Ҟh���9�)A��Ԋ��fs�a�8&LCCFp����~���3?v���kKS��0�c鮉�cs<����Z Xe��aa���
�_�*��; 9�+$�&���@�T ��+���A���qg��O-N|���^OZ�c���*�md�r!�Ϯy(��GS��Q#$�#�U/ۅȡx��J���ti�~��A|�(P�J�>��D8a���)��mG�D�/�!ą�*��1������* ��ڹ�;� ��9Z�Z��oN��_J���H�_�������1e�V���*{���)3�y*݉J;��������ǔ3��d��@���3�i�S�&�U�ڲv
x#��~���������>��s�u�Q6�!�?j�H���wpX����ᘪX���F��<
�^;�E+_ސ�6zx���r��Aۯ�w�`4 ��VV��2�0tۅ]��W�V1��лLO�B"ӱlC�P9���\?�:���6V�zwUy�TL�P���9��?rą�=?i�a��I*�HV"�5���������Gl_c\i�"���������}_����%�P�&C�s>�R'3��ƉU�o��E��qN��f.����X�$�Ta��r��\@�
`��*C��l �ؒ��ܬ�$N<������G�ҽ�d\��0���|x��Xb�]b��#��Gp�����1|wL��.�@Nrov}W�	�p�~ɳ�₝?���pb� ��3hl���]<��`�)����������٨�HTZ�Qd�x��=�ӛKT\R4t��&�8]�Z�T�?[V��+�_n����r��&��7�KH>߶��:yߖ�ғ�h�V�.��q>�����dt�6�+���5�m��D����FZW��INR�$�!_�kr��fH�wA5h�B�� "���fx�f��(�1�7Q<�$i���}r�ٚ��]��נa�"{%GM�ɉ7�����O|W!��3H��
8�"�
����������nQ���8��6.�l�Y���#�p[��IloS��1��>ԉe��y�m��L_�q/=���	��1B
3��vA�Լ����^�T��m@�:��uB�Sԯz��I�i����%V_I7��m����䐭��;t���aV��`@q��KR����q+,)�����2�Y5�3���~G���t�W2����-���J� @u��\*6�X��s��g���Ӹ�j�ᾏ'F:I�r�S>j��k׳�ã,s�#��"V��\~B\"�=��z~�>!K��FS0���t����yIV��)����M�U��-���&�
��<���&$�^dI@�&l��E�c8U��@�l�o��B�94�PO���p����5�%u����z���g���ؗ}u��R������!~v�a����8�߫�"�D�~e���A��O`>�s�[x�:��k,�B�M����M�����j���W����=r��M����B��V�{���H��2c��ƫ[��;G�%�>��3&���Ȱ[��҉��h
�j�!�~Rh��A73E�b�.��%���ԏ\Ԉ�D+��vƄ؇v@P�-�PǄ��Z|���Oz��7��)ݍ��<{�ց���H9�u��;6��(��?�f��;��W��@{���t���� phd�JiB]��,0J�K��7&ag���Nkzt�.K�0!�8���,�hm%��'d|��Y�G����3f�!m���餑3{�a�B誮�N�ޑ�!䨥���ٜy4n�mK�ϟpֹ=w�O�ꛨ��."����OP�"(̈́�Ñ�攕 C��>�zB׾��Y|=�C���h8XE	h�Ѿ�8�����\�[�3B���C��V�P&�V��&)?��k[?8Fu���h���	��i`ן�ڦw�6�o�-�L�l@�%UT�O�sDo�	�t�}���V)br1vAx1��Ҝ�Xݒٸ9UYb�u�j�k&�-�s��t���ͻ���w8Qu�F�9���P�Oe��#b�ו�M��3}���QCMbl

}��ڗZg)�2�r��0�N�I7V*��(��p�o���};���6&*V��m�H���'��$������%��C�TS]dZZv:J��"SL3�32uNl4#'�6��bJ�����
��}�F�y_r�����Mr�>���X4�±��gbyF��j
�8 4r�ث+[�V��j�S�����7И�l�U@��[YYHqtId��
EM v�
Y��A���������]�0�;�H�s�
�x��q��x�����j�-c�{��l�F|ma��`	NE��dӶk0�z]�`�Z���I����H��n�˸��N���1�Ee�� 8�Mm�F}�;��n㴋BDPi�=G�ڇ����ܫ���g���7x� BY�v�c��_��հ<������:$�p�^����ؿ�Gu(�� )<����{���E�Z�zPxvt�1���Y����jJ�d5�ngEKFpe�I��Gw-@)e�{&m7d�� �}��%���P�5-���3�A��%OF�DDd%�������p��x_���C9KB�
V�8��u��ޔ[{��?8���-����Z���y@N��e�!Oz�QTY�e���+�Da	�̦l�s+����V�"X�6E�GM/�Ի�U���jg`�Lw0L{��f��Ƕݦ����.�B�qܣ��AΌ�lE^k�5	eR�1ѹ�(3i�W�9
K�܂���˘~�_,\��NA�b�JH���V�/�sף��gY_��=�����;Y�I�I]T�==TdX������Z�9���2��?���Z���g��ĉ|�����)$�u;�H���őm���o*�Y0������`��W(����sd��[��'�m�)�M���(���Ss�0m7����Y�e���2��L�P��ȯ'�"f[l���������2AN1�}賹�^��`�&� ��Pm�Ż����е��Q����m������gں��zGok��3�n~��ة�Z��]��3>]�*�-@�D��פnIٜ�_�t��`��&�f8�=�>��פ����Z�O�YBgs�gc∎:��haih5��P�o��W, �x��ڊ�&�Du�M+ni��7��T���`��+�i�:9<��H�!m�z�g��Tr�Kخ8���'-x�y�=��v�x�*���Ԡ��*��hc!����`��M�f0c�oy.x�~C����I�H��^��q���N�2�[�*DT�r΀w(�	~9�#g�膧X&��x���h�؇�B�c6i�z�O�#��v�� �w�r�W�1��Wؒ�F���T���?���nC�5�� �� �)���.J_.��{ߕ�qS�[P�f���dn�eY��iC����^9�T�`�i� �@"�)�u/FT�|�����AWj���I_0�?<�6/�n�g+̉����?с��gG����}pٜes�7~ 8�`�����kN�����n��у7˸��ːqا5�giB�A{p4��Cf����V[@�5"���I�Wp]�������*L�c�9`7�9��[�ё�׶B{y�G6(�s�tؐA-�Y���EWpX�UV��xpS�c�4�g���K���d��h5C�٦댍	�|U����;�q�kg���N��d��Հ�S�=S���"�؜o�{S��r<*,uJm�*A����"`9m�����Z�g�ZǛ�U����ԅҜ��M�ǅ_�'���.Brx�������o�=�E��!�e:���jጬ���\����^�����շ]�ݵ����Jg��b���S�> ��D�S,��"�����酝��nVm����H���?[��ԘYKO�w_�{����OZ�7�� �m�[]�$WW�E,[)h�]�=c�Ivg�H��D|��탪i1�H�e��@�X32pX����'�@�xن#�9�&�YD�I�^�]݉��Bj1\{L�7·��4��,�X�2$q~���Oc������{�z�oܬ��>���>��;3�	W�2)��Kl��>8#E���Xy��R�r"m���cKD��iA���@?��P^�|�fW���<�	��(���w���߁�����0�<��:[��>��"�I�V���� P%��|��6y6dV
=1|���o�\S�7óV�U���Z���Q���ծ=������qam(��u�9I�����W�Є�~X�&#� R�i9��8�b��
�Q�'g3/GnHؑB�~^Z�T�{��´����Rr?��C�h�HU�r��A5�3�9��Um�t��������MF3A�q�C�pP�x��W+���F��n�%��;Zc-��V��I�(�F�醖�W��K<�!��ꯩ������٫n��"h�v�ln�T���WaОJR�C���Ⱥ�C��W�W�R��)js�F��D��q��V|���D���v�����ҝE�ls#"��*���fz�#�#1֙��k��F{��R�3h�������-(ڊ^��������[�yaO_��_�o�#,�� {$_�H���m�|�H�Yɒ�M��	l�,��S�&0G�N����)��
��՝1 �-k2|��n���������1P<5���V����V)��p\c���W�laː�Q$ܕM10P���8&u�$�NzE�$����8[+Z����3��`��%-��K�N`!���  ���T��
|S�+Q�����-׷^Y�Q�;���.v���}������U�m.rt�q��u+�j���c]l��jq*�ij��
��k��Z��6��,��:�����՝��d��LA����ű�Q�l�_��c��{c�ST��֪1�z�M%�9zF0�P3�A#�.l�]DsI�6��@�h*\�ଇ���+� ��g�u��J|l���jz�a@�X�Aۭ�ms�K��A������[�JV'����Cyc�@*��Ů��mȩ[�,�F����'����3S�9�@}]�+���W"��f(��(ȓ�+�6$����8`mzݽ��.cy���Y
Z��T��^Cۼ�.��Wl%R'�cI��l�'�ҩ��Q��9c�w4�]�^_%���t\��{d�r��rv��q:�ߛ� �<����?tc��;�n.�rɰ��zJ����_�k�{�5���a��h(<&��.�v���Y����~Qׂu&��`����p����<��1^�{P�,�O��DL�r5p���u�����:���(�c��N�d�R��@�o�pZ���d�k �2�d�R�KU����1���S��w?&A���aQ���XIkƉ���3-�;��!��8,�3;q�$$�^��aǁ܂6N!O�ёc�ͮ��Q髆[2��~��4��fZ�i��e$+v��+/"�Few�w�}��׊��e���io��ӂ�ؘ�c�ϓ�p�x�A��oܽp�xy�j#�z���_Қڢ����U�Mn@r�C�KV	�U:j
S�C1�dUȋ4 ���u��� IpS�g:����3R�ѳ��}�8����F�_z���z�����N6	r�\;p7i��d��[��Z
���:�MIL�����5B��D{��g��Mلk�a02��@.��=^F�bcb��s3�Sŵ悼5MEN��TQ�i��Μ3�qA��m[�\���g��z� �ϟV�<��t�$!�|�:�~��_��u��\�����)_���P��	y���>�Xs�&�5�n�2*���l��:����:Yhג�?��.6��T��;gC��B*}�x��L����.��{�F:���Q	��G���X%��pw�5Kn�\-�>��\*_���IA�^���p\�W�P���y@��y��ʽ�h8Q8`��$CV!)On ��G����Jrk�M����'^�M\�����@�Y���מ컽�Z˖ĳ3_*�հYއ�������Kڧb����V^vE:��$i�$�;���9�p�@�-��×%���EQ>6��$�Wl�W�'�9�M�a�y��"�M8�Fzr�O�zϰ@,vL>_�p�;��Ѥr�ǀ.z����3	�x��$����Dh�u�>.�
��+���2^����6G5#��'���p�Ғ�&�}��v��]b>�!��w�Ȍ[ct�,��Xâg�����=6�z&�ϔ����ᝯ��@�����2k�Ϧ�Z�+����v܆�C��Jdv����m�^�U����(dR*�Z�E��INO��`�C���O&��^�ƼbTF�ulWC�(�~��֠��;����7���M	�K��J}{>r)�רj�q��M<�ăD�����o1����E��N&��o�b�?^EN��S�f��"-f�(|Ê��9Ȫ�;.���2k����3`&C���}��?F	�'��cK�'Z��`�ɟ��7��ʤ�
��Xŗ&�Ȭ��Ч��=2'/��Π�L�a���2��޲yE��@|�ˎ�ؓp_)�����5�S��|��z��$� O2���l�ƅ�������7�^��A��/��8G9���d��u�?���y���1��hD~�ߏiyY�9&Y3,kGC�vy,~Ã��d�+"p��5�d�Ă�ת���Ep�?����kX�5�A{��Km���0�c���[�-PQ=LN���M�-,iD7H�qv�*����R�.m�B���!�o�+�1+��{��kvF�V�o��~�z�N? �"�8��#� ���"��K�E��@m��������f�e�e�I��/�?,�؆������1!��Bg߮��k�v�I��)C:%c��dY2<�gq��Ա���5�%����c�������.rՊ^�!!ˢ~����{�:�d���
w�\����f���f��zg�:7��B�"���&̺}��*o��b�@jbt�^rMYIx�G��Y(��F�����/�#��*�NxE!�ǜ7 N��M�_���<�!���*x�M@��϶����;3A=�b�����M��q����i:���qH��S�lU	�C�곸���|<�j)Q�*�ȿ�л&���a'	k7A��f?�O#��[�7������|��J5���O�v��a�wߙ�C�`�6�iό2�;Z�L�v�q�Q���o
n����?9���fz�C�u��D4��_��Ɠ�+��JH64��qؒGـ`�Şk{�
}�V�Y�Ā1��K��Z���_0r�M��q��z}�=�f�С.3is�ϛ�TVT�Zi�����e��=�Jp���u�q�F�oC׳M����8�yi��9l�!J���A]���%�n_*�8M�p*��ɑ�-�l�X9��,c�b�� ^Ц�be�����k���Q��3B\a�FD���_E�.���J�!͞�o�bg�_5����O��sEƙ<�x�s����o��צ֣n�/���Kɷ�/�*�D�Jd!> 8N���s_�hՓ����N�S�1M�)$�H`�S�X�.y�6O}A��OŤ6�� W��-ׄq��^��S��i*իv�:�,G�8M؟q�F��yov�"��:�6��&7�3kX���i����Su	��Un��nG�yC�'�]?˥�Ϝ)M� �Z�[�|��?N�"��B������a0>�M�A�.��Vr�^Ʉ�/Y����֑L����#��]�%�dW3�w���TFh�42����^�-���e��n���B�T��s  MV�%���������l��{��=�x��|2��p2���x��K�H���(W7g������q^T��Ʉ���69������!��E��d��b�E;��D�T��X�*�
v�d�>1��y���^��9ˤ���U_ZO��^�f�^�H����U�Mz�C4�F�E_��ue��HAV�&����S�a�2�S6��a���w��k}x�ܝ��E�5�!�
�pIjuHL�,�5��$E^R��t	�=+�/I���݄���3U"獟��Z�R���G�C�=|Ά��q*#��$��T�9�[��O�ZY��� �k�`pP�;����2����G}������H�[y�ė����E�tD�UD�C
{�M�
��Gֿ��޳.��a�{��W��Fi�Vy�{����ޘ���Ԇ�(�`*���m�H.z	F���]z`hW߱>��X���~����˝M��z��Ï��k��iq��ş�S]��O8�s��є�v�ˊJ(�︔3�9~��1��� ���5��k��V�5���0zJU	�����4�t|��q;Kb�bW��TN��$��E�����c�Cc�c��/��t�� C��c�!��;����sP�Y�dSJD��YJ�^��?(J�s���� ��cB�b>�ۣ�>��U�" U��k:.�z�N׈���� �H��() F�Ҏƹ]����_���{/V�[�]���(:�{��ڡ�X�h>u�ha�V�5��ZT	�-�@b�xЀ�:��lA'3�(� P����Ve�p�	�#x�j�c�I�h� �-Gw�h�]x�1��;�^l�Y�S��_��M��I_`ᐪ Ú�At	����F�?��d��9z����0�$�H�(��X�o$y�#�;�~d�4i�UN(�	ʮ�Y��	f�2���_���R���a��j
0`v=m0GB�s�lQ��^f�lj�΂7E!1p�#���%�i�[n<��4��t���tQG���h�i#�y8������F�Cj��x%�hѶF������Y����m(Z��`��n��5�(��Q�%[�Nb/�A�=ݞ�w�X�9�,�P>�"q�0��9�Ɗ�$��gq�km�~d�F�m�\6�!LP��0�K�#�[l�S���5>L�=��mqO:��ix��G�E��${�6�Ѵ480����E�c�Ҡ�<A˒V۫h�� ����{i�;�j��[�ѧ�����F������kr�r�'T4�Wb����/T�;���~ڄ���� ������o���G/���6�����a�v 
�gs9��K����ڦ�%5���ceh.FxA��ܯ��\;�na[i��wD�,��B�����|�GKW	��JR���^�1�e��?tv�'.���z�Ҫv�a:��\�oy� %���Z�E��V �����ٷT�C��G���uӡ�)�<�W�.݃��^�/	���D�No[
R��d��{��"kgA�C6u�B���n�R&4��9�}yG�n�tf�e��#�u�r�Y�L�D�EB`ϹS��A]W;v�`fy:��Lj!�dX��Rco.q��m�4Ͱi���jj��e����%�T�>���,u��V~+�����4X�@i�s=ɌMۆh��]���ÒC!E���������v\y"�*������r����v-�k��K���,�M+�FR�C� �RM�����S�����*{h��m����C��ķ��U��6�ZP��S��ż�,�J|�*��J(���m�ʂ���m��Yp��?�u�=��6$� ]��]AR�|���[��߅��ᤀ�qhD*�6x�ܦ�Kъ���U��#���N���L]�	\^h�EX	%,;~����!��H����ؖʤ�x
������#d�a����o�[���&$����"�q`Yu�4O�$�����@�/H]�&�Ѕ�몥ɲըߏ���)�����*l�7���$�;����gu��s��`9(HDv�[�����9�Ǌ�z�"��A�V�5�H��"6[�_c��,��V5��s�rI�#�������U��N&	Pj��[y3�8��5ͳ�kH
������W�����G�7%�b)��o�Sxe�-e�T˝oĴ���w��4�ԺG.�z���ˬp�����,��^Ŷ�8U��ިj��=�ߘZ.Ys[���;��)�%���4 a"n$����$vߗ���ao����i��%���!�܉��a+`��3��>G.m�J�0v�LwA��I�S��WE�9�:@�O6���?��\ŵ ��|���7ٛ��u�nO�1�H3-_��I�^2�� AT섴
j��	JZy���ܑ>�&�Bf�TBc ��� �s�+�nE��5�X3����-`w��d��Pؚq�Ns\NN�����vX�J[#�ݶ�`tDڟm�����(��Xzw����8`W� ��=+g�uo�vj�g�y$d
������4�O�?�Ҳp�ʎ�ݒ�V��^K۹g�'~�RFl�"��q�>�I�d�d��f<��9�q��+��IKU4R�}1��G�%b�	k�˽�D�U��ы�W���a+�n;���r���ݯT���(^��7�)���VjJ��ȷ(U�R�ΉW��Hڹ�fwΊy�@s#r�^��bC'�6_��XhПp�1�#ވ$\���R��b�������Z���e$��<H�:ƍi����s���1w�%�D���8�Ϻ�/�N� B���G�����[jv��B�gVW�C�鱓V٢�ܷ��Y(��a�b�9��i�G	s��2�z k��ك�	;�6��i*��)�Q��%�G�ć�U�	G#eV#�x��(Y�K`�gW_%B|Ջ���J���8K�۬Xf쮣����U㘊�
�� ���U^;�����`/��V�-˧���"���dG�8�Ͱ]̤KL��:?!�&��nM=yKyO�ۛ`�\�q��г��Sbb��H`CL
�'P�oͰ+Hx)h�X����5v�o=�]XM��#۸(Ym�ov�&ƺ���/O�I�iAF�e�N|�X1��!"ߘ������w��}�?����Cy�(�m睪��uA�]rvOj��pާ;e����uu���ËI��QD�$7&��$r4}h���x��	�6E���( hsS��9���9b��ѨF���pl{ܗ|�_��r�%�H����xҔք���T�b �>�c�����L��P����"?��e�5��#
1�T)�8a�_��J�<4�6��P�gl=��k��ll)P��f3 (��73��>�*����;�x/��~��ٛ�
j�����HqN�Ѓx�}�]���������b�J~�7��W�x��2�q�y6����p˵J�[��z�Aߣ�PW��FN�@'f�S��R+P�'�l>h�D��5����`b��P�3�y֖8��j#/�{�)h锺��.������2}vG��ꙇ�W�<ϒ�E����)-�e��Ԍ�n<.Ē�4�7/'��Uܬ?�l�B������Η���(T�Y�Qa�?�HŁ���1�9 _��U#����soA;i�Б6At^��<ǧY�k�u�4g6���-S�������53!/o����p!ʱ��<�����X�H*W2��ƆPy	B�.��g`����{�����*���p�*+m6MDV�M��@���IM�k���9�t.��)�Q��������P��F\����q%ce\2��|�q�Œ�(���ί��^��8A�O�*��EBrR�O�3/Eg\�o��� 3��ѩ�>��Y�Q[+�MM-���))VW*�5p�H���1v�Q���!��Z��0���06�Ʉ��S�Vem�A��Fv�eU�@���K�%m��Zq��9�qALr���|�[:nFy����D���YCz�G�+n�x��U�Y�
z�E���RI��EC�����kC�#΢�����)�H�
f�/�1���@w��^�.y|r�UL7��c����k%��^���ph6r��8�F^u͹8f�*�(��bt�ݾr�,�]�k8P�(��:�g�w��[ˌ(�Ej��16q�e�5@�hPl�Z�vQ���GMm��;�'��g�N?�`�^I���z��5���O������d�Pz	�"������e7�eݡ!m�N{�n�*�M�|� &?��.����K�m^(:g{MCRh>5ђ��o�Ӽ-�)��A��{���hL���\����ּ��+��[�Зً�������.����?4h\���H�}W�ՔxOܧ�dL/)�\D��&~�,/g[g�} n@�D���gD!j�eGhvq��(N=���G=���GV�?��f��ֳ>��m��� ��8�p����x��@�ә���I�ޑWGJ���/YD�A�O��8' ���Ս���Ԙ���T����%d��J!�8�zB��|J㪀����7��:�d�g�}�>k�n�R��{.�&��D��J*��HC��]c9����߈�W�O�0��-
!	���X�%Z�Y@�%k�mV��Q�A�bo#D��Jg�� 񿧯CUmE�O����"��\
�N\(652���*�}�)��3���Þ+�"��s=�I�D� �7�O�vZ�ć�mQ+���l��
 Qt���:��V]�E�ss��.��l#��V)��5�:�=x����~B�^��<	^d���üc*����W�h�Rw0J��k(�Ss.y��;���=�n	"lh���,�'�z�iQ�r�<$ ��v�4��8!5]"߉�T},����M	'��@�.tEf����Ş�|�_��6:gRj�n5�ȿ�������|K:�C������4}��)�d5��˵4����`<�զF^g���3�B��[,�h�����g��<4q�ə%(�璈i�2�o�tT�SM<��%	�!Y�1֩�U��1��|(����n��˅PP�-��#A�Sho�'�3��[�{'x�#��Ã��+�d�|9nr����2`5��H1qzLHĳ�)��5�c�����BF���ړ�G�֝�_������bN"6�c��w���bJ��}�TKK�:��|��:��>�2d,Q4�{Η�ڒ(H^��!�����9�;�i*8p�FN�����J��+�ֻ�{����kl1!r-Ӡ�uj�<:$���&\�rC�&�k�_݅'�T�����{����I�EĪ��Rٝ!v@��\�Rq �d2ߑ�֡��R|����I�ۜ�md��4�v�nX8�3���^��&��Hu�V8#�sF�}�����b7�[ǯ]E�E#�� �� � [�<�§�s���)����HT`o:�6�X�!�����n�~��	ѢW6�C���>;�^��LX-*�(u˅{�p���%V��|�h�H���0� -�ˈ���W�v^%a��B� ��PԐ�!�j�&�8���č�K�f�ҷ���.stoC���>gtc�'/�����ɉO	3N僆L�{�ou�iAh��'�<���x�O��6�;H'e�c�v%��L�mVÁU�1�h���wB���
���x�|l�8.�rζ�`��X�hG>Wn�m��7�+��҇��b@rB��[?�凕\��cZ���[�ZL�H��c�.oxr͞-|��~�?K��y��	Z���L��¡n�j�G��^u�B2����SZo�34?؈MX�1F�˶u�īN��\��ʉ��� �6��Х~g��R�F`�(C4�^�>���K#AM�2�� ��>�o��#y@�%�v�:�3�dM^�#/d,-��YĪ#�`Jos�F&��R��.;ß��ߋ���h�$d+_�-C��c�-#���@�s�R���/q�f$:�Q��
�����c�#5��UFs`�?�A�=ѣ��a1�����-r0u �t�K�����Ƥ��ăk��������|�ֽ= m���\��J��f�69|?lǹ�q�os4��Y���ɤ���\}�����yۆ�UT~���5�d`& �M-(�*�b�u��+yAu��ĵAlJ����]���o�L{|��?2mv�����z�t���yC���`���l���=��c>)�h8E>�k>upBRq���/Y'a���$�Y}K(i����mt,�X�4�h?
�6K�����X�~4+O������$��x�����<�~��9D��hК��f�;�����@<�ߵ�D/�!e���:zF&o�=��TG�,�)�|�vYL#h�&�`�W���Q�_rё��}��@N�+�;Ia��G�������"�7H�_{�����ئu�Dk��cVv
&+�˪�L���hr��ڜT7V3��L<>�f$
6c�y��`L�G���_+훖u�m�F�_���Q�k�{i����s1����6��͖ͥ}�]��瀬���D�s�
LMaI���	��9�'+��寱c�	Г�H6(��=㠻�"��~�+��e?0�ВM�=�gX����7��<������z�yFv�.�i��iɶGV�B3}Ϟ!�2ɳw1���a�3�[���6Җ�+�V���J�r���aN����|� ���Bʻ�2J0�32�tɕg
ot�v�b��
��AFD���/r�&ғn����pe�`�ήH�px���Q^���lV$����	�'*0����'P
�6��Y���$#�cv�T)4>����K��8<����;Bj�k�a@ࣄ1����J��/6f! �1�(My�?�\�_"���YJ;�ݵ�Hg�V���_���Cj�	�?-��dE�*��lk4����T�����Gkt��N!@������cdS��	il�uN�Jͨ��w}q�wM��fU����8�B1m���������V⺄Y���j��t��T�-���G�\�֋��9� ��ToG�������7�%Ȉ���l��n��6IZѤ�Q��,>9!�j���4��B�L�$� ��5��g �ǰ�L��d���$PpW �һw���� �}J���>Ř)�~g��)���	�U[-�R��?	�)ѷl�0#�+��9w��ĖZ��p.�e6�����/+��Wp�{��mO+k�<x�*�p��c�L�#�$�Z��u�'���^7�Ix�I�y����aQ"t��J(��?G-tr��X�"������;	�+��U���x�<�C��ox���I�U��gd-� ���e��2|P��*EO�jfw��������م"��#�pIT�E#�L"�:$���~�e�I"z.��i������"H�M[ aDԡ�Dg���Ά�_�$��V+k�g���m�wŇAB�B�����l�#D��p���RX���a˛ �W���)/�@@oj�ayۓ-ԯ����z��7(�Es'^�s/��w+�3NL�)%�흁��Yi!䏼6a:c$3$�i	�4g�q)�E����^� ����h:S'�5�U�q�e�|���d���(�^K5�N�GC�ǝ	���j�W�Pq"��O3!wc���-�����鑷�ƕ� ���5\�
%K�y�-�k��d�׊U�NP|��v���K+\���_+��>��]���G:F(�Y�BO5��u�n�)�z�����U�/�l�YU���r&Q!������N��u95�o|��v���e8�אO%�r��[ �>maX�ڵ�
�n2nl�+:�t�ڴ�ոm-8R]�Rǀ�������L�|�CZ�?.k�����5�ݶ#:Y�vJ�)$U����V��o)�J'�d��b��1��J��>Wo�,�O�w�P��a2���upG����R��zk�!�lo�C���Ԣ���C>�/ kx%QJ	���B@��5Dŧ���{��߿�C��:f8�M �V�d�ʦO?�X��y��Es]CU�R����*�,�0�GPW���@ˆt0:K���/���ob��C"�x)˦�lO�J�a�������-+�ٗQM������G�=�4�/��zv�k�� �j�s�9!���)C
6v*� 1(��uAHA�w�l2��)�J�{�_;4o�i�t[�du���lSC�6���R�r\���o"����JMa��X�Mh{DmD *2���{�F���޻:eg��[�[t#fyd^�ha�Șz@l�_���W�x�+���M�S���`A���l�3{a�����*�<����s�b04�(#�K�bGz�I.���[SI3{�q��p���zB�nΒ���Ԭ>s5���Gm�89�VN:���7_���3oq\���n�hJ��%�r�hi�h揗M�T���ϖ�o�C"��`��9%t����<����ؓ�ı���z��4q�9��;��ȉ��Ǡjx�/-��H�����&���WQ�7DJ�-#g���jy|����~����CQ�����:f�a�Ľ�\�N�KpÀ�\�oҶ�v�闹��C�R�z&R孈�o�ǜ��gPR�+�DkAp:�m���"��hҰ��B-զHE8b�����X�Zq�dh�	+Q�;T��Q<���䐇�#=�@�< <*[eh�����ȕ���R�\5\����+�ӆ��1�ĵs� �D�����%��vc2����A�j�!�H'�V�9�N�
�/�9�}����ނ��[�z�7��s��M��NJ�ԫ��̊T�<���,��#~���&`���v���<���f�����J�(�jj��p3����+�����X�.�����k%���L�j��n���]\
k�����5�+�8p=t��h�Z�g�o�	���8^�C�����x�R	K!�E,>�[��~����q:(�D��NN��[���{0%옌�S��?S,��t2ZD��5�ا��T�N�����`���&��m��!4r���5�˟�K Z�|�ꗎ��\g��#�
3������n��=���O5Ѹ�6qZ!����cI�#Ղ
� T���}�F$֢
��Pgao\��K��$��1�F�l��
=w�Gxw��n�T5��L��@a����f�)�� ���A�.�r���(6;
���Z.�$��|���u��uW�J��_��@be~��J�!��M�F7ג�Ɯ��*cU��!�Y�VC��"��	#����ZbE�z֙���F�?2�]� WXq�.31�0 �w7�½�=䷸����]�n�TBeG&���k:Z�8k�Bw��J�I�b@���2��I���o/x���v"�V/�.K5Qum��.#������^�+=���T_����X5[��h?\^��`B:��?A�j�{�*�������R�ax-�W��Y�5H�Ss�z����Ċ/��)G^�8[X*���Տ	>�1���)6���R�OB!y! f�惊��Z�n��	O����m�����` .=է�^ �7x4
�:����#�D�ol`pH�NfT�<��N{��G��F��U�̀�,&�u0��^o�aE��5�-�w]8�b�%貸��B4
�͢�bj����}`Ŧ�8�C+ё@��g.d.��n����C�J�����͟�r ��P18�+T����oK���})�}&
�s�,#|N(M\�c����LZ���c��_�:��B:$����������쀅�#�Ix��5-�]�Rq�Uܓ�|��wJ�6 �������49 �|�q���P��k�v-��0YQ�q�{���Z����wg���
�}�?�4Q+�����BQB��՞�WV�Д.t�q)s����hg�t�� �X��[�-��.�ќ����1�����E�[���>���l����ʿ|��Ȼ���;H� m��ϑD>TFz��@K��C7%"�b�&�h$0�����Q���X��v�-�}��Vu�G�;`9��SG�a�����������aL0j����b�	FI�4���rI�_��)�|�KI�JW����	ؐ���sv�7�}�I9�d �֪$%��./��z�.��uz欰26�ؖ=^�qa3E'a�`ܧ�'I,B��֪�\l��U�$V%hLW�;��9y3���+:Ӵ��gq)���k�+\RY��'����#� u�7H/@�8�)����F�㴨��P�V�=_��ZY_�.)�I���I�MW�������I�������)�d��t5B��|�Ey�8wE|�I�g��(�֟y�¢�W���&�x�T�f��g	;	�	W	4�4�\�ƒ-�R(R�?�eJ���[gT�S���h�$�V��)>���;�cߌBX��%�U��?hz�*m��q�A�ogT�B��m�&�#?��(�BN����W!W�\�!�8[n��-󣫾9�hm�S^Jb�2��\tU6l�U�$����&ֻ��g�t��1�pW�2���������zR�����2]xI\�,Ȋ�h�#pmEވ/�c���� ��|���A���w��-w� �{U��Υ�����}6����o� ��ijԶ��*�1��g
EM,�v@�x��G�5�P_���.��%<�M��kS*Ogj~���A�����������YP�0MtduT)n]&���*�"'����k�X�"\xK�zshb�:F�@�m�o���a���Z�5}a) ���X6֦ ��o�W-����<��C���A���>p��/�3��㰷���A;-.��L����-l8�f*�^SiO�8��c��#����>�J�f@aft�x��oӡ�r����(�C���i/�Y�/t�M#�Ѡp�蕘=���
�Q�̑���w����E#WIB�D0���EI@���G�?��v�"B�S�����~(&-�ڪT�Qp��t���_:r'A<�mR�]����pkV�ʫG������	� ,we�7�5{��*L����,���+^���s�o�n� $ ���B��Y�W�c���رq����S\rAVCZ3�m�n��#a�i|�b��6�C.$�`B�Q�F�{#_n<*�)�;%&�Zc����؅�^�3V�����R@M5���8�R0�dp4!ۢ3L��ǍZ�=��&pp�����2B���y��Ũ��5����8�=}�L�OE)�w���8W�A�'�`�$�O{*hb=]�x���@�IyS�j_M��;$l>�S*��]2���1s��%ZLnO�t}G"���@�5϶e��HޯF!��>l=/n�F9�z�ŵ�F���w$G�$�R�0�~U��&�N'��҃ݤ�q'rD�$fY�љM4�2�c��s�.8X1h��ox��X��@���u�Ѕ=O^�Z[��r6�G?��+9b)�l+���E�eʿ�h�g���
�M\�`�P�^�]� q?���
�_��/:Eے� ;s�����ssC�k��xK�pMc��ퟟ=B��SE�=e��0Om��:jړ�+	�<��s
��1g%��<�"�	D�tR%V�,<H{s�UY=�����8�z�������l����,�P�'��+����Y[5�Ng���F�����9��O�X�1#��P��&	ɦu'�V2,�h�@�x�fQĨ�ǜ�r�[d��#F�}3R%��!%W�g��\�p�.w��T�9~(z�ay��z�;�j�����G�_;�#������+*A�g�� a��'�6�Y�?;�d�'X��<B�H�
��
wD3Zi�Ǐ"ry+6u��?�p5_I��ɲ�tD
�J�a�|T��m��E�p-��.�R�b_A��\�z��]@�z��4|?���z���6���;�k�J
�(9�	'п�H�̬]���ً��dC.E�v�d���!�,�3U@�%su*�>��+��s5f��>��Ҽ��0���aY�2����Z}/�`�g�0���|�o�����BɈZa����YD�#�����''��#��)�1��и��t�\�BV�>���<�.[wqk�5�1K�����r��P(�Y}K�����DK�,��a.ѯ!͂��+ ��z�x�|Ⱬ)�e�UK�1YK�V�A���,(e ��8�mҜGkk!�_�+�ͺ���岂���0	̈́#��)E4�+z��hF�8@P{�	���#����)\���(Y���t�[:�{L��r�G �`������H	����>~"����/}u�mq	���a���,����`�n0��?�Ѹ������6"J�6GƲ�"f��kR�B�T��0~�(�P�Yt�V'�蕢Of^� HT��*�`�*9�2P�+��x��1�*�{^��R��$y�Q; �ւ����l�n![]<�.h���I�v����P
#hR��Je���#}�qh.I#���3"`�H�ٴ����q�1i��\+z�'Ґ��+
̔63�K��Ħ����XҲ�e����2m;@C�(\Άq��q��
�V��c���Љ-���)�NA���~C`�T��/���F� j�x��ǖ���f��8gĢ�>���(�}}�"&�8���A2�ﳹ�m�J1�w���9���&��}U����o4+We�"����%�	S�e�P\����xm�� =I6��*�0�A	!좂�,��V�l������v�Ձ9$j岫�%��2I/<��]y���S�.��yt��>�s�0'��H�>WsQ΀ct�e֡6�'��A���ێns0
8��6;�@�/e8_т�x�v��׵����(������K�������݋�o��A�D�䢬\�V����L��D��r��	.�A*}Y���+�� �	"�
�a�>`���݄��L�WOr`�؛�(�=��g�@�j��^f��pW�?N�i�Zu��2�U��Z���o�D���y}�ML.S�E7#�DR�4d������9��n��:�'^m�I��p�J���	�%~�G�Gz�1��jZ=ym�z�ڃ�'���aR
m�M:�·n�8X��^��{
���j~5Ϥ?4�קA��2��e���'�A�tL���;)\b���YH����DC��S6��6L[�$4 F�h��'6�A�v�)\x��oGܙ�-�c�*���>@0�D$5�ǝ�,�|{ uG���7v|^�O/{Isug�-6��|��IX��8 j�-��H!.`�����y��Ote��.Ŝ��{� J/��_۝_J�V�N�Oo|�$R��,�-�j�����<���$�Ēv����������C�$�)կK���Z�����m>0��k���W����[������N���~��Ar��Mר�i���GU	d�o��)pB(�	_J��Zae+��Ƥ���ṼB4.�K�V���=2._I���F���Y�{��(�3�v��T*)#�,��%h�<x�S~�Ԩ�����Uƥ���k/��� ������乲%�^��>7����C�,�]����1ݡ���[!|�l�4C���w�~�qpr��80�{Bi#E3��������T��Fte}��+E�p�BD�>��f���}Y*G@}'u+���Xb�*-_4�C�Ҡ�S@�����VWi7�b�i��b��|��x��ѕ7a�*Z�4�%�����I��T�&!�EH�+�QOJ�H$���2s���1o���$��ky<#Q>�yoH^QW!%�C��W�v'�s�Ǥ	Ϡ��=Y'�X��	�4睸|~1M��jh�[楻o-}��V��N��`R��9,��/{ɂ��<  D�=��"��I[�d�G��Sej߀��z�L�3̯�$�^�����WpZ�����u�o<<��R���͊6\�tp�d�f]��P���{�[u���B8��7"o	��ڿ���ŵ��Nknp>?�N�̇��R�d�3�o�k�T,��qz��s �57����ݖ�.@Ė�^�Y;�!�}��ä�v�j�4�v}L( ���zn�w�iG��Et��I�WY�Q��5�=���$
�H]a��7��Y�Yf3�Uɵy��˩��oP��=F 5B��-�3�oj�q'�*L�e��sFQ����Ap@qq��_+ !�vb��ʻ���<Q40EA|�l�_��Ф)|�Y��c��y'}@�}����DQc������D|�t�A=��˧�*�F��Գ��6�z6$�����VlF�C�~���ގU�����ץ�O� 1���E�ai�,w���ȝb�NZ�>�uoĸd_�p}@��_�!I�� 7��`d�I~�^�NF�D/�����on�>[<�
�9��P�@�L��	��90+�����	�2�	�5S��uO�f��Q�S�8�<6Z� R�E쌨H��*|��T�>��
���58Q�T��՛	
,w?�PrqX `k8���|�U�ȗ.�m<�C��%Q�ϒ$�l<ط9���iHH�ث8�ek&g@�V/�裷�Z�J���¢�k[��u�į4'��u��)N5�!%.�3MH�T��Z���k�/#�g��+Nk�a�Do-��}�W�9���Iӹ���W)��	��ȿ�I3N 0vYz�n�B?���q����<�o�Ż�L�r@>VtBv\(4t_���B���/��!�K��ӊ�/_��q��U��q��5�RR
'",��T/�ՙ�Z}�op;�4*;��5�{h�xm���%s���ag[b#U������C��iݟ�KFD���n�n~.�(H�����^�v2h������G�|8��n�x�b.� ��-5�_l����^c���@O���fȫ�7��;�x-�ֵ��jX|ܲ�B1Q��&@U�w�Ou�M�;�:��Z!��&(����iē��(�i���a�� '���hb��B�5�����Q���Ĭ{!�dLjEH��^����F��J�]�5�2�i���z��?t9D7���P8��N$us#4*3�����X��
q"Y��&�^��
#e{.:��żۗ�ʟJ�G�A�V�@Ǖ������B1�j)�+/γV�sKf�Go��H�ۖ���C.�PN�JU��,g�fO����h<���\����$��a�x��b]���X��r&��c�n�Kjw��0nZK�y݆Y�b����i}���H\ڑ�^��ث؉�:mz7ޟ�g'�I{Sd��),�E�Ei{d��L�N�3�-`�3(��jM|D�ͣTy�o �a-ޣi�jC�s����}���qKҟٌ��� x�Ȱ< ��Gj@u�
%��Ӌx�c� ~j�C}UT�`��4���9~bm�J�K�25ef�7�}~m�!�3N@�b��γ_}�Lh?Z����� �)�v {��IfI�cB/-��Ƭ�h�$ˤ�K��
��D�>�$��Oo�¼GΥh|�z%�"I��R�)E�/��GE f�;�>�I���+,u���|J��]q����d!�A:�������
��W����^�X;L4@D���6�Il�+�y����j�we�����>����Z��$3 t��	�'m��~�4�t(�6�,�[��!�B~�j���'��ӷ��t�E�"����å�|I��&�����e{����D�����)�2�Bf9�6{!wyKg�B0qX�b�%=�
�����
GeDx�'*�J��5P����Ӊ4�Z�ZQn)N�s��)�N1y*���z:8�e>浫g��S-we�[X��T�q@	N��9�Wt�JS����He- �r���7��&:Я���F.�F�bi]9T���Cah�:���@�~��	R��X�*�d����@�d|��{;�vV�g�� ��Fg�7���'c�����A^E%���e大�6��](u/@�/椙��H���#�"��Z�b���7�h�k�v��`��ƤhH,�!�^�`�|����3w�\ޛ���!e[���
BH#�"^G"rK�V��q�7�%0�M����F��~$�S6��?� ������{�{���4��ϩI47e5���QS�aU�9{rc�y�����^l��5۞	bmѻ���򞪿���&O�EiI���{����:�'��ݤ;���(�O�8Wu�i�u �H����ޘ�W��Ip�M���N?�
ͺ�/Jj����z�N��:�GZp�/�-=�֡η!g��0l���3 ���O�B�9��ݶ  &��7�-*y?�s�,����Nn�'n�������\�7X���ԓ��I��v���qf+"*��!>q�/�hH���Le.�`���jy����R�on�
5 {_�K8���>5&���XJ� .,wX��
�"�֥���
�BX�`���obC+@�9֋��9	��5Q[���ΤxTF�ͻ�6����� m1Z~کlaDc�>�މ.9��CQ�8`m��#�5��p�7�$s`n�3�|[xq6\�1�'� ����� ��e,/�-������ 2�M�ˌ����uG��+H�����4XB<"V��p�'Ó��F�[��,��5(��P�R1aq}����X�J�������<�Q�6/(ۄ��I}�F'7�y��{�mt�	In��>�Pji�n�I�7�T�?V���<I��E�����Z��C�OL�G�C�m@i�OFU�A��5�ؙ:�6��|c���[<��q��&�;���/&#F��P�a"��=���(6��ۮ�uV�w����D	�+��B����;� f�Y7k��b��4�C�z������B-K�x��� ��P� "��,xK��}兯��!{x���L�cB��9I�5Cv2�6��<��[������참��N!���FP�1��r�2�v�¡33Ֆ�-뼣Jx �|����8�}��*s뫻�Ɨ��V�e��,��Kdzc���C���.�p�*�숡FXH����Vk���ۣS�Ӽ2���wPX�_ż�,�[�W���|��
��f�O-i�HՂ(�Q���V��%���L�������4���A���r��k̮�|y����}�7��oI��>�8v���Xp5�\����\Ag�9��1��ϭ(~�����q�ᩖg;���׬�3�d��,=)v>�Z�9A����0@i@8SA�LW*�*�2��<�Bm�*�Rt⇫ԍ�o�r�ԩr�	2G��*��J��L:�+��G�ޅSB랊hD���WO��v���mLM�m�-�4��ߓM����}�D�W)����qd��!?W�f��U� :a��,Q�f�`U�;k�����/�E͇D �(;U���d~�nf���y#F����UJo��
C�P\����� A�R�_;l�y��N_
M�������=�RL"L�v1un�8���*#��Tߍ��<M:�\��]�ݾ��~��D�uf\*��;�S��ys��jd�Ix�]��i2�Z��X;, 6���`5\$Y�rp8�T�zC����  �F�Ti$�F���cJF���t�V�_�c#=�<	E�	����{�9� ����ba�C�ʅ�����W�pS\F�B\�)�e,���w]Ps�4�gO�D^�6��=>~�*�J��=+�Q����6�f�:h���:0cV��Bp�p[�!���F�*��ޥ�`��U�]kz�]�F��,֓Ag�"��St�ǧ�.�����1_:�,�����5�%�ᐅ�Oj
όd7�멪��oN]teR�M�*oL0�wy�c�qOc��
o����λy%}��b���mnU TQC�r<�������}��
���U߲�0N'�	|1ʞG*D�}����U1�J��2m��2�>J5����h��j�_\j�O2�GV,�K�-~f2�J�F��D��t�%Kpw/�I��g� n0D!Ú>��W!&�b��N�\�O�@^���<�Ց`�\V���zNB�o�K�a��irϣ(WÜ��:��G���y�#��A���>�{�m� ��:n)Z���ML�.`� ��i�F��w��:c���$�9�gy���ﬦ����{i����G��Jߊ�Mk.5�K�jM�����3�	3�g �s�x	?[��� )�^��n���k�8�٨�U}����:}׻;2��'�O�Gw����^T��ًhBN������[����G�Mz�r����>�}�zilJڒ���I4��օ����)��:�s�F��%0��p�X�7/��lzt� .>��J�s�v<6�ܪg�۳�G�1���U�B���t����� 03f%�CQ~���t��KA�ӹ9�0�,�-�>����6��H����5�Y������sa����q��)�����|�L�I�dV���dZ���Ma̴��x%�Z��x#�����t�gVFͦD�^�6 �*��-����02AR���{}�@��{��Q�%�#��yR��+/ 5�\�h����=ϸ���,�_}��.��/�Z�w��3%��$���]=��.��}m9�2�MV����r'O:G�E%_���M�6��"n��&�STD��͏8�����cm���E�">��qY�iN�LR���g�_�$�M�A�B��1�&x[P� �梭��IY/�g�rf��D���5����[�͸� 8��M.��tC#�������H{�˭r`�u��W�u.Bul��͉��wg�^ԡ��G�2'g��Mz��zP�ss閐���g�U1pɸ�����Z��}�ä�C'x��v�Zl�	���9!��7�Se�]�xU�b9�ϲ�/>d���̖�ٚ��K��Mwa�YM��^�$SG��%2�n�#�7�%�lS>a��)`_�)�)8��%��FI���L�L���i���]N��c �Ҧ��O��إwv�g��~`<�X��Q��X�.,�ȋ����Yт�h�I��m ������Q2��C*�<����V(d��#^Z�n�N[�f����A�)�B�����D���7��
��ǭ/u�%�,z��q��|�,>�I��V"���� ?��?�
�D+r�?�ܙ1�w��g
�m
�3��7�O�MV��ދ}i�4�
~r��]��-�?��g�O�g8���F���/���B����),��zJ"tj. �Ga���fl�Y>}U{ը�P���h�3��]����A�7��:U��w�����]�{'�� ����K��4n��9��ޔ������:G�� �J�<�����6��m*�JNbD��xr	,G!Ld]/�G
��)4
8`-�C�d�iT�nPt!�74t��)O��K�b�,�
6�zl�V㗪���ٗ�F���]-Hx}!��_�,B��fx��F*�Ap�^�K���!��Y��Ȅ}��Bg}JI��!�{N\HKO\����� �LUl��3O6�u��� ��r<ՐZ0Q�/����Vc�?�4�:q��6�,�[��~?��B'���g�ٯ���;F�G`�:m����-�����ss�j\-X�-o����v?�RL�<o�H����LAWfY�sD��ǉib3�0�*}Ak��d���cE&Ғ~mM�2ny.�ym����*+S�qY�H,f�u�l'�_ƞ���HS�;�ۓ���|Y���f��wd���Lw/��a�\1�$�,�%���C�NL�D��Ǽ��Мoٍ�c�ڝ��R�}�Zږ�JW����\����Ċy9��M�O�'X��
(�Zz"y&鉗I�_Ye~��|���OY`�T<a��Cʄ�|�I�bHO'� ��/4,� 8�D�l��O"I��z�}����V�dfG�h�G�yӐ���� ��y۔K�;�g��t^�5@�@i5d����4��չ��4�tː��k-r�Q1�N`�����o��3k��Jɬ&�=�k���v���錎��oaw��h$,7
���˥K�4]g�f"'"!��9'@T��2�v  ~��G*}���XpͅD�d�$�sO���4`�:�5��*�<�C�nݩ6Cfݝ���\K[�&=g@�����.�h����s�U'7���] �d��Łڈl��"�Qq�(���?��/���0+�%u�r�]ìRn����aL੠o�A��F�����0[�Y��������,�k�0Z���v��&�|	-ax�ɺzny���^9Ä1���a�I@75Ol�{�,��8L����l���Z�����:UaYw��j��]T-{�$��XM=���������?�}o��f��=!�tfE��Dnw��*T='�i����=�J{^�X��}(�y��HB�zz:���/��X���ĭ�2�[���R~�z�z�&�0�]Qm"3Ap$x�w~�Ie�@R�X�"��x�q��fH*� ���UӐ��V��I�p� .�����REzOn�w�0_�Iq�gV���u����~������݈����H��g�4p�6D�8�k�����+�:� �d�gJ��a/�S P�|��ǿ\s�ۄ�FW����1>��s����P\�k���wms�&]~M$�ؑ]�?v��^'6�t;��jl���>ӳÂ���@<�"�ٷnz�9�f� ϓ��6���o �8A�z���������V��3�6����6fn�,��^o �����	g���0N>3S���E���H�B�z��
�Ͼ��C��Dt�U��Ŏ A���͍���=!������ؑp���Q���ca���Js!�G�����7t�S0څ8n[�;������	b�8�U���PyhI5a@�C�z��<g��X.u�,�eҚ�%�ڈ-T}G�$Fa�(���[��e_��:��5q���räT�{�E�y����~i�Fy�T�!�K:a�%�����/����tz�M�����I�	�|�M�$E���A��$@��<�(�0�P�����јs�8Sdj2x��:h	�6�b����D9<iq��_���9��c�X�Ĥ�Gү�N�P�a�1$A6�"�]�X}���wJR(�l3�s5N!���. 4%!ʒ��v|8Z/m��2�}��7(%��8/N��=�
���}O���}es�P���Pr�[�u�ap�O�����pd,�2\���n�]���Ha���9��d!�J;V�����U��s�����	��&cvQ�?[�聈�L���V�ѓ�����+=�j����&���W�Sr�/B&Ga�/�1����nf�6�wa����L�x[�D�B*� �d_���^3�����Mk<����RDd̺����F>g5�j���	-��y��eb��a<���\�	��+=�v}��d<��K��m"ʰx;���8�$A�N`��3�Ρ1�M@p�%!ܩ��B*��{�`ؕJ��[�i�7�Y�������:�B��[f��;��I#���\ܳ��k�C$Mh/ �����޹�u���P�h��H��̺h��G͕�(��ݱm�=�b���cڂCP@�H�����G5Xxk3�$�/H2��BG	��J��	�{��Jo��]��u�~/��x�DO'¼B\�k�C~��s�9���g����@�2�$s�$ӪQ3��G�f6T��)F�ǲ��j���������a#��M�zd�����G׽���}�d�|'*l���=�)�
���"kP���&�v)����2 ��no�B�_����<����L�3y�Qǌ�W��RM����v�xv��EH�����v�kfN\�s3� %}���_�}@�ᨓޙ��i98b�UP�17�l���ÈNX���zE���bn�u�*(��R�a��u��,*��h��Σ�f��4Jp	>��L�x��9�t�>�⚱[k���W�6-Z���>��}���5+��2ܕ��	m����/9	�]f�4��bW�$yQ�G���QOw�������y�W� R@x�O����)%� �3�C��<$��q�̍AyR�5�6��t�8�?�W�{Y̷h� L��i���+M�`���m���f���5�C�Da�/�X�{�bx* =��	+_e���ZJf,X�=KAR!9�R��a+�(��h���kc�k�h'w��c#;&76�K6�;��1��ء�$߇�r�+�s�����`����:)5&᧋�$�6�>8����,����|H��]��ۏ|�]�,�pVo� 9.���Hgf���%RAqF������\,���4`1�Zr����b�7'����.h�r����8�R���b�ySw�"�U�)$��Ns'v�%�j�/H� =���U$)O�>��{�Z[#QGML��b{5^E�f1+{��y��&�$K�)ݜI�β��
��V��jtڮ5�"���ڌ�	�aT�n�j���:�Y��[�x�6�ڋ��8�LUgW�ګ�i5�/��Q32nRX)wa���x���t����E3�n�9s�)�E��~�B��E�����%�	M�)^��=�����1��pӊ��c�?�_#7$�ܩ�E�B��?詢�F���v�`_^<w��`r�{���v�Z:���^�+Źi� �>�1Rͅ�7�z�-}�� ��W��,�s�,~���H�����H�s{���Q5H��y�礀v��V]�s#��jѤ29	h��(Iqm�p[�.����oę�Bz�X5-�j�G|WJ+��~�d]��_�
��;�v�I^�=PՒ*��n0�an�8�u�90ZW�_��������0�_h.�Jd`�c�٤�\�_ո��]��KJ����J���O���ݻ��%��;Y)#J�<��Q��=S��¤[�l��j� x����VQ�z4����g;'(� >���|�GУ��X�}M�2�W\c�A��ƃc$Y��%dȕ���-�^>�_GN��a*�=B�jN�k�&�����v�=rT1B)��{���e����B;�^�B�Ĕ%v?�3�Ɓ�
�~��m���.C�b��O��a����[1ޅ#��X�yζ�@��������F�8����0����n����ğ�]z�9��Q��M���W/8A�G|Ԁ~6�A{ԵC92z<�X���d��Wwn�twیU����]�s#ۧ�}_7�f��fbq5��	7���V�]%�(TYr�����0s.��ytm�6���+�/�h�m{Iy�}���3QS�$R��ΪNY�:�c�b�Y7%Q���Zԕð=�W2�E��) l��{��bƨ �/ﳅ�|��Y�+��:�IEʥ��(I�d,����P�K�0��<�j�[���&�b��>��jÓ{��0��Q:�/�j��.��o+�ߋ����zQ4P�Y�R��i��<~������Ogs~W��G�)�U!|T��8B�w�e��(��˼E�jQ^�-�܂t�N�J!��A�%��O�˺���"��krʴ\ɫ)"K}�|����$�m�(�1n����s����Ȱ�l����DcS�	fP+WY�?09l��{l }�(�/����+JC�=гF�]�f�g�.�[�5����>Y�2|B$L^j�$+.j��!U��������h�v�$	��X�b�.��������U�B�:�}�&��!����>S�����	��T]��"�SQ��/Ɔed'��",�.�	��0s�$�f����D��>�Ny�ۓr�'�6"Y���#�1]�FRx[����+=<�1zת˭�5,���Þˠ�F*���8֠w�Zȷ�2�RT�X�̈��������b>�Z�׏�A�x�A���pLo!��o���x�g�Q���׼��H�qCm����?�����?��+8�+6��H�Þ���:5/O}ɕ�/L1j.��{�{��� �*7���3R)6|��dt4�c�c�>MOX6�c-^����:et�2�X�w㦌�3K%�* �c����׎���s=�b����O@/��
L����=�+є��)��|j�J.�Le�e,�*AJ����	LE$�P�� @�|<N9��|�"����¶�Q�2v$����vȚA��H_]b;�)Y�F�Mb�w��tYOW��L��W�Y��(}t1����'`�;5]d>�?)nEm����
��
�`������i����9�g�	�9�e�M�N͎�f?3�G.���OV�ܓ@� ��,�=8�^�,��	�V�u��t1��Բir6�Ùp�4:و����;�@\`6�k �9;��2�+�' �I�۹#~T��$ֹ
_��p_�B��2
��VfOf���&��7vx%D��xN�j�$X� �`�����K/�����"������33e�g�\�*O��)1��ge��2�'�u�z!L�Nq�\h`�C֫�)�:�tY�<�e��Z�_Q1rN�w��)�J�6�H���^����b�EW��W3��@��4&]���̲a�_N9���w*j����Fva�,A�F|DD:�:�OI}E�~;1��y�߂��>�3����TZ5��AB��j4���0�"iA�E{aT��ə)���ŀP�zpŷM�eξ��i1��|�gA�uY90~1������9��}F�(�!�6Yd�m֫v�����be��1i �ʺ+�j;($�r�Q�͕�H���Z�� !�o���J�'3����N���jKz��D(�rdJ�K��,�w�>�^���t+�.ǫ��>��NҠV��#��jw�M�Bº��Fi�c����c�� ��bw����vs���{ѓ^;��b�Ҍ���+_RސG* ���I˃ݬ��-���U��o���\�/��I8��}�}	An`n݉�{�(wx���.�³d(*k���e�$(|��Ʃ؞���w�M%�L��W�AS�Y�C3�:}-�w�!�@?�{�J|E��I���ƝcA$o!����!��;���@La�$��7��j��u�.
J��Y���|�9��Ɋ:Ec�r �� ı�)��s�k���6)�e�Mq�Ay{$�S�z�=3�`:�U��Z�;S�ȤV��~I$DOdz=�<�S.�1�H���F >R~�6�,�zb}�qo�f}|��ӾH��@ڗ���P,�	��X�����d�t�&�á�mnï���$G"��5N���ߡ�(�!�Ѭ�Z��=��s��S]�Wmte�XYuNRx�OS5�M9zn��ҕ��r�	��˷#�''�[�K ǀ��v%�4�-���gsC/mc�%�E����6��(��D��f�����v� r�U��>cZپ��D'�$��}�f�����Q:��k�&�8u�wE�h��
���ܓϏ����VZ�2-����a}G˙�v����A�LV.�	X�Z�КM
Sp���&�x�5��7\\��;��{��I�j<�zx�W�*Yך�^�B�l� 9�9R�"����pC��CR��O;&gg���0/�+�
�Q9\��ټLHu���=������6���7y!ə?;���{���r���yv���Q��ں��/��.��905y�|��J,Z,?/ei"J�n'ٹ�tpDsѶK�z�nxz��R�.�{GE��_i��Vr����'���Q�?����Ѯ�]�h��M��97(#��H��,�?s����@��:	�w��g�BW]�}g!����y0a#e���ٵ���!J�\��%��SMue�
�<��x�a3�ɬt}�Ur���pWJ�e9(� 8Pgr'���Ŭ�0*�.8w2�,��Y�]VNEG���Kl��Ѳ�)��!��ymqb���>�����<Ӎjw�~�qʧ�Z�$@.��[)���E�]�x�^�1�a�etR��k�l���N l�� ���c	�(��	��UMbf�Жb��IU�,4�t�]�x6&�5@�IÕ�Ӱ>tQ8*Ki�n0��{	��C'���G�|�����ͳe|^+����<̑�(�GɊ�gA	i�2u��To�L�$���D�bK�ɤu">&z��MŬ���g�dptm�&?�����R�֮��BUGr[�x�+��O��C���A!�8�a�8(+g+��9ɒ��/�8C�Q _!������#�)E�>�L�ѩ��H+N�E{՛=&Qr��B�N����[�ל.�sl
��������m�D�S����*V)�ah�;[ƏqG��	�,sn�@�})mN�W10��l)����щ�/�h���6�)��y���q#���Q��y	d,�|Vb'w>#�\�G^~J�+��[C�a^�����y�_OR�AhB�V����ٻ����I˸�Y\�w�X�%�#�/_���4�-w+��aL�p&.�[�!�.k��C�>�K�rk��-T����{�z�9s�IEL���W-$��BT�Xh,��h��<2h�#�YE��"/��B�>�����cu��p���a���:8��Ud�K�w?�&�KB���ب[$-~=��^��Ɖݒ"���L�FB����-��>�2=W����Z���V{'k����'%�!Iص�t�������~�ٷ���cS�C��}�ͅǳ:}u̹����LS�%aS�zTk����
6�א�HaG�3Rf�_��g,���Tm�w�Ğ�At���r��h��Ӳ��i� �h����{�^�I���2���Nkư�ņV?kWY����z�Y��(Y�}EO�g����(b{X��Sw��D�;�2!Q�s����`����s#;؃(#��M��N��c�r�S>�V�mbx;<��Q��x�W9�.����$���Wz[�Z+Ӝ�3Z�[�'h�-�כ�뼟Xk<U�>��x�$����S)[�i���h.�r-�:Qy���=ɾ��ˤ9��Y����$��ӧܗ�U�~Ы�~r���it�Z�ҺZ�s�<tBpwO%�����{B��$����B��Ajl����S���>�_-/Ԏ� ��]��S���[_���p%�<���<5��r2����Q�L�����Z!z�i��>)�;�[6��Ů�[���'�S[�{X[��b\� V�Ņ{U�wK�{b>���(��~��6d�~/��|�1����/�wH4��^_,ݯ���H.�;M 7)������D��K�X�K�h"F��߈dc��x��D�����a�~��y+i��+�����b��x{r���|d�2,�>��V%t��Q}�(%����rE�?�1�C��5��'s%�IK{�ƍ�wk1�"��뒚��1�<1�;:a����8�NJzp(��KOR���_��j|�i��H8�-���=�j::m/%/�S�ܯL�J9sg��"���=����W��-O��o�-sxW/H���]B �6�eV�u��Ȕ��s�G5�&���1f�
 <qN#t��}�Ld�A�h��G/����M�Z����?�X֭�6� A�1w����eG�f�O�蒿$BZK"�����y���č0�7s�b��kp�n��W�|�8Y���$ﲉ������$vId��^�����ܫ{v��Q��f�#���`���!��3a�w�JRx+*�:���0�	R����gwneY���YX���ٵo�� k�v���Y�7�N��Z�צy1&j��:c�V4�׆�_��RZr+:nIRC�˃�YY�f��"�/*���Ι�`ܝ�xi��L�ҤX���L�q��GƼ��H����.��]�GL��i�LA��*���ⶹ�A��O���8w-��%	Sel���>8�}�g��+��DR���F�a������i�nbwԌ�5
����pv5�؊�|S(G²D�%�������&#��3���ɟ�9I��Ԯ]���U��7j�/hs�OIt�z�t-⮡k��Cm1��OM��
P�W��=P���g!�O[h�~}�?�(���ݙ��g��uw���vM����+�~�)�s�
5EuN3��n�G��f��C�����ݐyB1�>��,f�;�Zn4y��3�u��N���e�2�ψ�S�N%��^��{Ȫu;f��t��V$Y9��Rm҄�-^WC
�U$�a&���\h��k�%o�:VɋW67L}�M��A�!�<1�S����9�w�-��){~f,�}�!Y��rY�/�Zp�ff�3��ږXM��<�&G �"�K��
q�8������dX �I(��Q1U�\e#�ǅdH1|�c�||�|od��1�`�V�����A��(����G�O*-�I ������e[�^(��S���a�ӎǕ6�dv��	M�l���V;}o��l6�3����i%��1ֵ�ag	�� �c�o:8��ӕ�eJ_P:V��up����a Dks�Cr[��ݕ�zV�B?�RwzYv#���%ֳ$b�I�K��>	��d�x�F�o���L��#�<�!�怵�����5�ާ�02[�t���v��ݼ���@E9�Є�������P|��=1P0q��-	^���mG��>�6OD'q�� �XXZa|ʽr%y�O�4��w��t���:DG�(�ʃf63������� �����Y��aY%�Y��m�
jo�xw	�<�]�9V��l�2�ӡt�g�y=Sʨ]�g�v4�Ws0���W�@(}�p���H��/t���V�]�~��h%�O (���E���M�$U�I�eh�Ӑ�͡-�� ��j8��
r<�Rs�#̻vj�Ğ��2��W7Y>;���H)$68���*��Klu�&0�u���
1���۸;������q���m߁̒zm���V	�ťٍ��ܣ�8T��*w�CHA)¯~8���P��_��h�����׮F��c��V�5���Ψӫ����Ë��&g�W�P�r9����+AMd �!���SݍoMLN�զ2�ђD�0�.�U|rX�D��׍�ye���z!g�'E�4��'|L<�l���e�{P�	OdԹ�^�� T�8��i��h3� wr}��U��3� �3������9���^F�#G^���F��9�l+K/���fܵΦ�M<ʕ���ׁ2�
��T�)�)���wZw�uxj�b�g�d�P&�G{��ϵ!�p).t�9֥{{�į؆����U�U ?� p d�K[጑��ƽ�j��uu�@G([�� �?��ߓni��^�x`�H�_�"Q��o���ל9Q��}y>� ��د��3�m	�ҏ�-f5H�bU�-�\�Lg;�km|�߸�	�>�V��{,,'��*VY�bjT��U�W�����I���|�P��
���i���~�U�ek�)'ֺ�ۃ��|���s���V���T�@��/�����iԱ��hnFPւ��OB�ͷ��zK��S����8�!��_�Y��9�z�ʴ U�sK���>
���g-���'C����)}���70F_bgfQ��1�&M�}�Ke��zF�s��eه	��a�����	���&� ��.w4��oUՙ.y����k�˲��a���M����C3)8ff�뚿E�u:u�tH�<,nK���u9�7�4<��B�j�ŗ�mx:15B�ӟ��7����s��0w!2>8��Ş2H �A�g) �ݱ=�ŗ�;qJr|\�s<RϝPh,[K��y�z��w�sރ�����aJ��SGcs5;f�o0y7��q��|����'w�̀�F�D�%�U�%�a�����=@��Dέ�? �9��kBI�4����74n|b&�n
-�_��BD{R�'L��3T��)Zi����&j����u��<�Ƅ�鬃?���-���_�O�~�R$���u �bBɊ"�ðײݗ�\�mn �1�H+��E3���{M��$t����ǚ }`�Z�{�N��y�o����kKO�7a�;g�X�6V��_��,˔.�x���%�8�b��T�]˾��dhÔbj�s-JQ��|F\4"���ʷ6 �ë�����>��w�y��_�L���#W9U��˩�$O<��u�3�;�ێ���}9|t�v��m�ßA��A���.�T��|��ed�_uQJ��c꺅���l���j���+}���jY�gz����n�Y���d��˘�9�z!"&�o�����p'88�i}IG��}�5�� �IZmb���(^���"2�}��C�Bw��`�p���"�� B��TƓi����J�{���h�C�?���,7�*i�> x��(�,?�1�V�}�ʡ�M�q�D!�53<�4�'�Y*
.�-3�2������S�=�I��I�p�_�<�'�4=���06)��:4�i����_�-���K����4�&�9�x��܎���������=֤ �����4gN1�4�
%�K�F��U��ӏ��{5��@�D�f�F�em�nD�Z���s5|}���Av{�nF����<�XJ�����w�3!d�6-����������Z	�ր�HB�Phk���|��K�|*��?nY:*!ߥ�{�����p�ܯ6��=���l�aȠ���
�=�:Q��"�U���dZpx#�g���I�x���fx/����R=A2�z��jA構s>Mc�"�d�j��ET�0�zeC��9C�g��-߂���,iT_-s��eIC-2��`���р[^;�i5�=\�S{Ĵ3��W�,�ȿT������^������?�L](pe)Ʃݏ��ҢuL���5�9�q�;���Qщ� S�'����Kȏ�p�wi�&%���8���ޱ�Ӟ(@�n�q�6�ɝq��1  ��B�f@`l�j��.c���������qb��ec�{�?��LZ��̔/�ö4q����{�v��noj��N�.$5a��[ZZD��1n��K;�Yͦ޼��}��;�+iy���;�"����bN*�?-c<�zz���б�s o��e2}7�s��^����m���Z@%'���iu�ܸ�F�A*E��U�9�ڊ�K��W"[7��G���9�<��L�����d�������l�.�Ozk�)��ƅb�R��Ϫ�+R���t��ŧG�l|/P��]���Rɩ�ك?��/+�Ȉ|�n\!�[~st�f\y�ߣ�zh��)v��B���ro��sL��u�g��;A�DH\p�9xu�X�g+a����!��tL�NWPJNaR'����R�/yQ�$�O%7�*/-�1�Uf����b�t�C��<�z�ٗ ��������&�d�lO��ڇ���5�Eti��e�xS���Wƕ*��Vհ=y�.^\���|��'.�| ���y�'˄�7�_L�;a9v��<��G	]���?��=V��f#
�u)�=��M��G0��g��j9;D�=;�	����V��T����9!��=k��M��8S���aT8G�S]��||��Vᒃv�/�(�e!2#�f�p�\��0Ϸ� � M�B�k���q��g>�a��D�`���uQ��",�PTo4z���4�T��Jj5��XQրtI����w�t#M�hV
&�:�s{�踚�V�z�g�K'�;�)�Z�g���[�[aZL���R�s6m�j�ڔ0���l޼j��8�$��Ri$C��.Okqt�� /��J��
u��)�q�EI퍵�2�h>[B�����沋��)��D"b^���X�IΨ P���L�^�T���c��+}Qtdj4����f2J���/#�a�MY��u��94�
�X��������P�G��2�U�����;��GdǺ���U�g�f���c��;J�ѷ��ܕ݃oܬ0�Gjl d�|����
f�l�9��!e0A�M�<"޺Ӻ;�r� "�{�q������`6s�Y۠o<<�T9F37Hw���8e�ve���ikF�q���U���ֵ9���}�L{���M��,�6%��$��r��hܰ�B�?t)F�ؐ6��4�;Х�t5�����93����z��EeIߨiS��p�n�ҫ�+[7�>�R@w�D�?��f���G��0A�[����Ֆ�/e8pe&!��_��^6.F��F��ؼ-���[��,W�HE��(w��J0�������K?��@^0|oF�l�&���I]6���y���X�Y��Ux��P:�v���qg F��I.�hu)�FS%,��m�_�ʴv�#���Y�?����K�j�H]&��m���j�p��f�?��/�9� �樾�MĞ��\-��^�ݼ�n�9�DK�������3	�E����&��OY�\�F�B�05�a�%0�U`���[�hǊK�~��,KK�q$��d��n�e��qF�9C��������t���e0q��3�\�.�:��M�n�p�5GvϠ�ͯa�SMd3v���'B�|*���y��	��]l]4e�:�g�0ȷm����D�zQ)<C��5��8g]f�HT�?��:]�ʼJ�P��]�L�������� �a�nK<���1)��;�9/�ugG���;@8�y�+.K����ĜI�L
�a-��;�+
Z#��JZܻ6��Θ��׹��Pe�������PCZ+F�1�q�j6z	��ʐHk�PJY��8�	�d�o�h�\���nM�v�["��G��j\��䐏ݭ��D�aM�I�bJ_�_�Jy[
"o�Aؖ��{�Ӊ9r�@Y' a�W%�_����g<G
hˏ����!��ܥ��lIu�b+�Ԍ�%��8�ȧ��Oc#��a�nC��e�T,�r�(��u�o�e�	���cQ ~�j�gd�B�1�v�^c����~��\�5�P۫&��g�<�?Gb*�Q�*�L��F0^Li/H�Z�����Rܛ�)����f�� \ aK�%Io�.����+�7��j.��3�)<�>�1|U�!��2�"�O��I��_ ��c�^"7�r���
7_1�V��!��A�|��*�]��t6G��S�|����8�P���cD�}�F�ه}]a�Ґ8<�m���z5��A@�9 w:U��w['�k?�z;��t�1����t)s�L�U��i��q����Z�+E?�f�{𖙚�N�|5s�#M�7dz��0g�B-Z(�,��_"�&7��G#/-���t�R�K�'����H3���ڳ�L��/ꗀS6����$�Qm�8�o5n�������D���ʰi=�j ��c�c�B7K�]Ļh\C0�.���J�NK�'�� ��^_��A�Ǒ�w��c}� ��ϰ�G��*m%�EI>�`����0]�~j�����+�J��Ui�,a��.\�eC�����RZ��@{�l���|���
�j؛��L��<d�`�b	5�������p9��Y�p����������e{���?S��?.�/ �4�5���ŕ6��J�16���E9���3�]�2~��d������ث�/����n
�4>��� "�z�}D�1Q4h۬���D��L�,m��u�T`�[�1�dz�0YH�f߂M�k����:^�!	Zr��RP+�5/�]���xǃ>ގk�j�ӖC����\X2n�,Z1��e`	�q�(Vm���$H�$X��J-�e�f
v>4(��Gp~�ٰ����UۈRۑ.�:�T�i~fV7���h�D��I�i3�w�i�z�v���1��C|�$��E�K��k ?�DM��Yܻ�9�3�t�����LТ[��ot��9�l����e�
h�Q��k��p�^E]��n����^�2W3G����PC���I��JK^o]\v#�q��z�N�X=6�ѣ�5���6��R	��z �|ɾMKj�xqZ�5J�ͅ���J����o�l�p?��N��9��V��K��-r͙D,}�_�e���K�Vxc�]�:�<@��	-�H�Jܭ�_Ԋ�*Z��O8�v�KU���:d�z�M0�Q�+�lr�{&H���6�2`"J�N0�L��8�9>�;�r\L2n�s�B��<��+�ߐ�s�*:�U���i��qC[L�}�]fxo|Ɇ �Xԧ~�zB_�UN���ND�;�͌^N	L���	�h�V��fq�ҍ1�C��D���l��&�H��~d{l�6�$;�8���̹�͂Z�J���<�nC����b�8;����@���]�����>į���j)�U�:�b��+v�4~b�,o�By5��_�"�
�6C>�rѪ
��吆�4�@䥴��
����A�P�a�m���Z��`���k*]-�B�VH�`M)ЃG~�1�w��25�(U��6I4��jVhy�!�6�k¹��a�K�\�o��C�H�?����c�G7��͆�g��9NU�\�V]��f�̒#�-�������,��d�RD���I��r'頻G���	F�7 ���������bS�_��H�\����_w_ ���L'-u������D:Q��l�2+����!Z�P�V*fg^V	A�ѥwZZ��{7 �����#��^�3�K�S�GM9��7��-�N�u��7�w��f'5u~�=��fX�\��E��6����~cv?hH�Ey!t>[��:��6/N��ю���ePb+o�c&A^� zo8��JN46H^	L�1��ma�[���<�v;�^Zw�_G�vq�X�nw8��ZaOF�`f�W�����7]���P*��VS%�'`hN����U԰==��P56tL{�]B�a�%Hf�#W������${�?��OOF+�L7Z���>'@qǇ"�kӪ�;)�s폍h�Z5��	�25ц�̦�+�\���Ez�G3�Ŕ�o{J��Qk2���ń�հТiU=�V�SZ�E�h0��s�v��
?_q���(� �����Z)��t��PL�7KL�� ��QA��w��ᚒ�i�c[�-Z��w�"D���g*���Va֏�)$�Z!��C ]��ӜY��h�%����߽��� �7�R4��@�=~=����t���:���@�4�
��%һnP!ۃQ+�
'��ki�Z{�m��gP��8!���Oi	�:��~[O����G6Jy�Lg͐������=���R�����h�n��:.�ɨ���6��g3�����դQ�W�2~��	�%RHP�SIhZjj��V|hp�z���SQ$�sh;�����k m�H�C����M4��c�!�"8� �|xs�AGDS�'���W��W��SaĴ���P}�Q�%,�F���5���t��*~�^S��;���k���֞vUQ�U����4�,V�>�K���Br+��Ȫ͔�Q_z��k#��vJX��c�ʐ0��~t���]5l���`Bʼr��F#��8}�1��>H���n��S#��eK��SJ�t���>X���]��/���Q^�h��e8$L��T81Xϱ�v��A�����o�dR�L;��!V���^�8X��	�U��v�̤Mq��S&��ޛ�)�Xإ�Ԅ'wP�(�ci}v�xNwaQE�Z>I
#����p�t�{5������d~0���r�Q(���o$)_+s�_�5���|�Ǽ�o�Hb��:/ڢ�U�O�aY,���L2b�'���E�2�U4�ּ�6� ]��i��e��(
<���|�ZN�"f�b�(�A�}9Z!4�8��DZO��ĥ<��<\l7F���Z�e�x��!�c瞌�u��:�o_G�A$��f�
:��E��ъ�+}Uè��w,��
^잣��F�ב@9Swэ1S�g���~`� &���lnL{΅���$4K�0�����y�iPW�%$��2��
��Ȯ�#|S�j����uuK�yS"מf F�W��Q��3㶰״��(�B��Ҿ��$X[��{���>sҝ��Z6��t«��[�x�U��*�Zߊ�^���]���47}5|~<�C��/���96KE���+K��p�\l�[[S"���F/ZS1�����}�X>@>�Ǔ;\�������$��� 9fD<V���x&֚�<w|.6�t��:�S3w��Y���\ĳ��{���}�A(?��&*vqz,J�o�y�=�o>�@e{�6^����l�:�%�0$�A��ؕF����ftL��{�ȗ�4k�~^�ڤ��
�&4C:r
�-��@���"��`Km@Z\�к�5<31'@��A1�K��a���U�z�ܾƈC�5L�>в��
�T�&�k��)�.�K\B��PWʥ���=׃�!��R������*�C����������	k�
����h:2ew�k"��~O"��������l���<F>��fLU]^�U� [��z�G�I&eV14��<}�Ӊ��G��2�{�0�D'Cr%t����iƪs�!�¡ء���9f�rq�i���w���K������zp��vt|�.v��TN�գ�����)���e�i���Y��嶘6|��#�Jo-)��l��)r*�|���\�Ap���s�[!��L�i�V1G��M�\܂&����2քQzx���&�l���l8i$�~��bE�֖2�w�@,�1�Bϊ�w�6���n�>{����x��M:����C���*�U<�7�[������	�X�7zO��^�i �w���I��"�O������y
�;�����scu��6T'|Eq$Z>yw�A@���N]i U������lR�����:�`����.�W��z
n��.�ǧ�:~fh%/����"�#��(G+�lV�Yҡ�E�� �0��l{��n��,$~��G­m�����V��i4�����f�Ζ��'��n
����y�� ��`�$��a��`^��v�vǏ,�{u�I���Y=�kq���"7�d������p���B�D��ZJ+�"��Y�d��2��݈��(E{�s�|����%q��f|6~�T�cX($��6uǭ�O���*9���*��]��q!�1���,R����j�YD��8ޘ@e�	$,���N���ȵB9��u���RBb�}X��9
��WT�Q,��4�"�[J򣸻=t����#�²�������h*�#Ƥ)�,�������v1��~7��ji݊�E��X*�S�us���C��T�5�J��������8c^�ԴYs�S���c�s<����G���lځt���o�a��-@l�ӵ�\h��,#��;�8��F4��0Ld�x��[a��6sp&������;�l��9�7��	�e���ZK�w����J��q�䎹:sU~�Ch����m�]��v�sY��\�q��r�|O��G e2Y�`7�dN��/�?�:���ty����^�4��	T���Ks��H	g��Йk�!�z���M>m��N��R�7�򪈵� �x�8�+��/��pϑڡ����L����'��fy����4��K���1q�5�3M�X�Z��ycΉ-�MA�<�>gh���T��\�����!�[��~Xߵ%��B�����K��p�Y��hI���wuV�c6�v��|�=�a�s�Y�q���F��Ķc]q(�D�,�.n���Љ�����&T��H^ٳ} ��/<Uä�IV��	���h��=��_1P�&�<-r�C��<�3Ԏ������f}E�Cn�M�]�qXt���ZN�f�rdd(V���Q��z.W�=
/�vҘe��&��Ƭ	�2��Q��� �1���L��p3�Q���^z�����c��.��8>���"��ԅ2#ō(�r3	'�]��cΩ�o;$C:���ե>�0q�}�pStI����֕���?ҽ9��9ʽ���`P�����4��w��
gb��tы]H���H`>�d����:ڨݠ���m*����M[�{l4Eh������(G�G�{:��/��ZZ"̀�V�c�-e5r������<CtZ����7��C�?7����2=�네5^�����b�̡�M�:��� �Π ɷ�;WM{oX�PaO�?�Q����?�R(��mIA�'��O6t��6��9*Xߴ�����`�[X���m�n��B%�2�/�(�$�F�~�H��Vf�+V�wNzw�b��|H%���ғ(�f��r˂t��k���4�d�V�����f?9�\X,us������6�LdLZ�?9#��� ��I �H��	oj���P��/�m���(��O��&=�aU��&U[����6�Fa$֔w�Z-F	�؁��U���h��PĐ��z��h.�Xʧ��7 ��D|1G��x���K;�S
���� bh̝4�w�Pː��GT��f[M+nvJ��en������;���w��A6�	��Tߑ�'N��Y��7:��b��3����Aw��?�EJ�/`��WX"\��CL׍�w�<Z/�8�w"�T,�X��`���,;*`A�^KM����QKuU6Z���S~_;��=d�����v�17�߹5�]�}�I�v���cz�"�Y<�'�gߒ�Ò0� <����a��e���>�N�����Չ6�p�>geL�I��ypr8��9n�3u=�Ġ%@�u�� ���m�N��t��E1q|����	��w���#�����n�.������,�6'4ɶ�d���?�d���k/��=�a>��^���E-б�n	_�ї��35J�N�E��I�-T�~�K�j���/��DT��v�Ě�>NH4-�g����/۲t��+�oģy��[s���K������tRlSS�H��U�������k4�S��1�kyE��ȣJY��m},��5v�ݎ�!��d�b�c�ICi�
[V�u��_�i��o���3 &X�	'� R1�W<8$�W�+ !_���}@.��+|VR�x����F&9�d�R,��x�G^�Z�n�}�hFwah��ήm�8le��&��q��zX�8�" ��3�cLN0m��ByX��٘��"�ޢC�u����R��4��������}��+4���J��D��U���qy�t��Y6lQ�6���ۇs�o����C�,�H.W+��`�!����">��>����`j�#��3�Z�B2�z��Wl���H��X�tR_j�̀�EDb����V����$��?�gzx^c��M�!��|�G�Ů�s6L�W�Ea �D�qARA��o8���@`t�UN� �E�	�K�b+�"F�we�}��T�zhe�X�(���0�~x�K�=S�7R�לh�k��Y�`���1V'���3�NA}�X�ڴG,~%Y��gvZ������|��bп��}��֍��W�e�P��8]r
����.��2'���)���[�9�ٝ�{}����B�f2u��)H���>�����8{(H��d��lD�r��<kB7�<�3xe�+����m�~Y���N6��͚,�aw2�`zD���҈Z#L4��{�>Bq�Wv��f�n�U0��#Ɛ�"@�����Pr���|���@�lb�q������y+' I��$�������A	�7T����F
��{W��j�����=�z�R�*E��HET��ޕL�)�J�,�=8^lH�6��:R��w+L�0��+oR=�̺��TC?w����d{��	�آ���8��g����YJ1�s6��|��FaZ�+#𴰇�ĉGL��������DC�x���VF�"��K�,^N�L�0��Ȍ��ڞ�	��\�o��m6}��+����'�-X\�R���3|\m0���� �ʹ�v��!]�z'�����-99]5�M��������v�05{�u�ũ�D���O��Y >�^F�G*ж|�s4<���ܡ��Z�sJ���c�� �/%�V����CHU,�;�EÍ15%U��)�Mړ�k�3���[��x�V���m�{]��K����=?���B\GF8��w���4G2xy;T��*�c��q�~b�e�����hgnV*�NN�������E?Wp��Ʀ���<�S�s��F"�V�F:"���Xd�W퓓{���[:�A��|��?���߼�:��|B��K\�&]�
�N`� �8��<�y
�燚�ŗ5z������1f�W��r��$��]�����[���gp����r��:(B�j��Ҙ-P��90L>�D��m�6��$���!��>�H�P�!9&��Z������%3����~�9+�W���K�_���Ou�W|y1�)�3o���A���=��ח8�1q#aIhƷ��A�u�D����M�ˊ�'ȱ�l�ޣ��i����}r��b��8w���Ԅuj�%�&:)�]�f���Oh#H���T�	C&q��{�K���:~wr��$+�����%TZ�(��K'x\�cT��n<i�6C��]d���j�㷰�m!����q�gDui����������H�ú��*}vTI�O�&z��`��OFN~��2�dku��yG�ƟF���� iu�s�.i�j��ι0�Tn�� ��i�q[�?�̤D1��vX�H�Pv��5���W�q���]�����l��H�M{�����N��ў�ۍ{Q��ċ��5 ����сU
J��9 �MR�!@;�ԝ�N(�<��[�����Jn�M�fb�X&�m��L��a!�De��Q�����Q^j(sM� ]��Byx+tR5'z�?�R�|�L��k���plw�	�Gyb�D�誻�>g宁��Q�}¡T|�:��Y}�"�W�.C_k����չ2h���eUd��c��"ԁU-?���Mb�f��4��y`b]�*X1˻+��~F�2)�|E��#Qw��#m�/mԆ���Op��	H�Sl\�$2��6��\�w�|S���8���y�pL h���v���u��#����8�F�kQ��FJ����s���F��8�C��E�mj��/��f�j�0�t�����cd���T
�"llԱ_��%���&RC�:�pb�7ޚ�?�����h����w�נ8��I�ґ��Ռ�nK!����2���?B� S�~�v� @��� ���D��]w0�z7٥�
����38�ó��(�m6��H�ފ��(?x
ù����*��Wi�:o�>�k�n{PP{��X�RFzI�ߏ`���Y�d�Y���~��%f�u�ꗕ�^.*�ĖG�������,`1���(ȀY��O�ԩ��A��U��^h�@�ri�Ő��>	ո�p���|t��G�"� �f� d�6)��k8G��F�g�|.���-���Qm�/�v��W/�*��&W��Z+N���'�
�e�h- �t���3���}���+��k�zՂ���X|4R��b�i�xe|J�׾C�.$Ϧ2_���-^?LBj���*�F���y~]n��̕y����R���L��@��O<x��/�͋+^E�.�*7vk�������q��W'}�$ �c���������}]��޿K��K���$ ~Q�[����ï.F��Snn;^��p�hG��s��9�����}�:�Y���'�	{���mP�r��-'� I���`��%����rg�ץ�־��^lq��%�[Rt�̝AѬu�Qx�6���L34�$�c��A�1���D���*�$ h��+x~�>0w�_<��C��S�\�%NՔT�}��<�8���ob<�(m%<�G�1�+U�����k+:̅�B�ٽ^=�`�+����0�����+L�|-�M߁��p��'x�Z!O�o��Éoh����lĺY4ۧ�b��	�5�xJ�{��c�"���Au������j#�v��P���D�:Z/ 6-�P�n�c�+j=�Jh\i�D��ߦ���%��z3/�&B�}�<��F!��2��V��̽�+���i�'7�}gC/+sc��b�j��׃�ٞQߚ>�����w����[(�'�i�>�kY���zR��L�S��������P7)�(�gut��b��f��0�� �^��h�]6����pN�r�p�4����r��/�%V�ږ��l�`RR�*X j�i�òt�˺Y��I��wo��Z�ØK��&�i����%� �x���=�ʿ�Ɲ%�\�x/�(�օ8��[5%�e�x���H7�HA��U�=u���a�8�n*��ޖ
L*���0a�9�z��Ҵ2�Ƙ�	���c<���3�O��q3�<�k����7����Wr��Ņ|�U��"S�N�>�a�������ݶ;'���~`!�IU�0��,�h0dݳb��y�Ҍz$ ��ׅbEŝ�Po]]��%��(%ڎ�y����1o�S�Sdq��1}�*�<�7'��@�%�f�Ͻ���ʰ5Hqi	�k��*����f�A�s�M�H���2^��Ԫ����`���h(���˥�4��a���G�.N�CW~����"�e�L�8,�&wd#k�M�3�3����m��3(��ܼd������!�$ڙ�<���,I�C�Y�\�>�iEK�>��,��.%48/ Bj���<�;qo�	��!(־�K����T��!�8�Lް�Am��n��r���[Jlm��i`,�ۯ�tF��
�c��2CG�iz�_����.��@p�W��
l	#Vp�n<z�f;ܫXe�����=튘����Mk:LR2w)$\��+��[_�7�U��5����*L���`��q]��c�r��f4Pszx_������S�h1��,�Mߜ�'X�l����cz:�J,��1�]O�Y[SI�C�q�����s	O�~}��L.�[\8�0����w<�RoJK}�!�� d�W�9�WM���_k�kUo�a -B��ލS���sHܿӫ=!iyu�T2I_VJ��:�������h�����M�&�+�W���󌚺��|�x{m�ϫ��˨��gnh+��I7�p�}��3�*�\[���Y�+2�O�i#V|Ss�/�&��\n(�=s;���d�؝ޛx�!_�>�zԔ2�99�Ӛ�0#����T�}���a����SI����"1�}��B̏nz$u[�]�&ic� hhΎMQM�����qd�G�ա��ջ�ȼ�ɭ�Ϝ���4�4ފu�|���v��M@=�3��*𷏂�ѯ�0H��%	 KT����Zn��n����a@�Ϗ���:3��`�%��}Li�|X���J�w���X�)�ȋ�	8x
�i\e�G�]�T�7(�U7��"��y(�m����2�hf��0"���[�.9}��/i KJ��Eb�����FGn��T�5�H�-��B?��1�S���@��ЇI��s	~g���0�S$7;}]���S�nu����F{Tϣ�}�\�p��)����~�����hpn���Vr����`�K_d��%�S$	�/�}ֈ|��a+��Œs
���>����	ϣ��MQ�@!�����4��S�Z�-�Z��r���[��'N����S�F5��?�6�bd�ǖ�5��b�:%����"ً)����/�н��r�B��B�/*S6�ޘh,��вH26pfk�֫�W������{m�s������q�F�դ*� !b����7i.�Ʌ�y������a r�S���9s��*���j�vl@$u@ ��=j�+�MM�DO���-ε������d-ڪ�J��攍R���kN���&�L;@uO��m��g���\��F���2���5��U�Ƕ�[ x�����@��9o���@�g��6 )�":>�����I�侞�XQd�o�4��1ɑ��29�KŮr�Z<��=��>�A�D��"wZL@,_"5�#0��'��x�9[�N~� Lt�vR;��on�5Z�XN�:v�Ԟ��|h����FPfz����MXKQ��o �ٿ�ǘRy��MK�0����JD��Qr�+�u�)�PMSU�i~<�t���X��S٘r�� ��
������s�Ԥ��ZxE�@f�)�#o��.��-O"�)��.E��+��:�o�\��au�nя@E-
�A�R���k?pR!���A̩-Q�$ރG*�g�U=.�L���ܠB��R"��Ж����gPI�??�?�ع3򕃌�U�3�H���(5��'�.I�ɨVX͈}�F�~��FVL��'�]�N����p�m�v����ɳ\m!F=Х�[ʭ�E7��g �E���������:�'�$1.�����8���1,���)���gYc�F8@��a��m79'���^6���>�)Pﲲ���b�`��tJ4�IbYpGTt� t���K5�"ĺ}D�/R`Q��9���s��h|��:��	t7*�5X�u��djfv#�0YN����<�@�T#z{a*eR�d����u��b@�,��ᴱ",{���l�u�8Wc �E��2s���P!R�P�`$�&�n94�
�f�~��xI%�5�?�k�'������5�����Q���^�
����{Ȁ�l|��(Cj�:<��k�nB�Q.l�����@{q;�wڒ@�\:w^M8$�e��$�X��X0W�.֫���t�J����kP]:E��-���:mȡ���cߓ�����?�)�o�&��L:�T'@��T\��2�V�h~�W�0�"�c�Ԓu�y%<9&�����BiAa�j�qZ�3��T]�Q%���h/Xiw%H� {g��Ε/+8;�,��#�����z�c���?;H~�����+��sy��|�:). �Bۡ,?�؈�i*?3U��*����,�������*Ji梷��1*.�� ���8PZRQw�+XH|
W��H�H�U��T�?���`c@}Z���R���!�ۊMB�_��3C��P�Z����jL��+��J ��x�wrt=�g�0�?���=�f���3� L%��-m���N���zB�랉\)qݪp���׏��4�k��qQ����J�Y*��|�^'ZY�Ф�ZRθ3�%��J(������4�1J;���Q�0��C,(M;�;3���Л.?I��W�� VG��ɛY|���		D��#`'c�����4�y�����7q���ܸ���#�s���(��u�-.����|*�2���6� �F�T� .~'<��N�]i)M�(�1�Wyѥ�b0Ė3���C�۪�4��Pn���qh����[��c˟?';E�<�����[��Y���Ӟ�j�(���Ay�Y�� ����!�]��[����ֱn��b�� �8�/���Ϛc(�v#����~���@jF6G�:��uo˯��	ģO�`p��14R�����bD��N:�B&&b9��#�q��H�`�L�V�6��f"��-�J�=�%�-�Җ��yb��U���3_��?7��f݊��cеI7�� �����&��%�F�N�~���#��q�I!@�+���
�FE���-���P,bY�Yhkՙ����䙜Tg �$�V.�i(f5d������V|?Z�c�OU{\�ę~*2�~U��< ��>��G���EV��0�@�N�4����*�=���B����Olw� �A������g�B��ˊ���{@-n�]�r�ۯ�!�6G��������m���u�Pgd�)���/4	����cHk&�CER̂��=�i}J�Ʋ��]�j'_ �}4�����y�u�e�uOTY~�:��J��Ks�$T+#�;�(���5z�a�%��a״�f�c7��Ҹ��9�hf���4w汜�1*)[�Ϋr��}n����z��lã��\vN#K��1J�fK�ϓ�Gk�"��,�:zp�_�T�۱���S��l%#��Dˍ��3Bu]�X8���T=I�������06�/�b��3���Z��Fu�@������-�׾���vE7yO�!,3
���.��^�!�:�}��g�)^�pĚ�j��pN�{"�y�4D��0Ǝ4Z�-^7��!PU�^�f@��j�P˶�,���Cm���H �k���s���/s�����޳~���3H�x�%a*����9;��?�<YuT���!�K� �����(ɰL�\���	w�_����(��s�M�_�$_fD�|^��/�҂���'ؐ)�fo,y�^P�|�bZ���Bm������� �u��p�0_؉��o����qe�K����Z����F9�y��ic4�s��,��):e�8�oeZ��.��"9ߟUOU�x����]�&���F��^�ZO�~H��˻����oP��j���9�b
 ���"hg���^k�|G�%B �����KO�.S��0.��z��6�`aF����h�ïb/R)o3#�}�O{�������"K�e^�"o�ĩi6m�J@ܒ@"������&�~��������s��z(97���QU����o1փ��h�P6�R#�����-��+����≞�b����9P��г]M6[�7J���}�yBfVGD�O�(�#.8�⹂��t4�R	�lN�2�a��DV��v�K4_��d ����x�	�O�݉�12�)��!�P���d֗�K{-o���J��@�s��*���"K^����/.�'���U�]�w�#2W�l����0����dGфK)�*/�����]�~t8�ƕ�t7�F	�,���4�$�v�:�#;�r~ZA�c6����g�
���u�dS�����[��%bEʒ��t!1�u'>�����^']�s�4T��m�K�I��ʧ������M��"D��\Ѩ4�Y"�W����^4�uk2���D����P�r���\Mi����έ��P3p����OEj�;1H|,���*����J����L��c�{��{h��=��]��B5�%7�!o��\ �ct��	G�=&u�FQ�t��[��(��}ѐ�r0@~[J�G�+�!��l]����9��ֲ`��9	�c� j�?��h���gf���y�Ma�1�Ldk��t�=�.'�p���&�n�C���#�e��;��Jq�?i�ͦqԢ^7��:�Ay&=[ܡu0=7�PYc��`S�c�3q˿Bj�x���(�+��ݔ����)��ǀHPm��&N�a�|����y���F�����v0<�`� �h���k���ε]y^�(h.?.tJ�	,FE��Đ:�s�W`��i�ڷ9'���0���-n��3i�ְ��%NpO6lR�s��ާ��6nw!��lO�N��V�X:>�$4w�Y~���N#���#�y&���4�H�j��ьX�8I=5mִ�`��y��N<6�+x�C��5���Xel ���Gt[��0�|�:��K�6<�t�\h$��%#�:E���2-ꔤ���Ŝ �/	�J��������ș�}py���?�B*D�2G�/� ?
t���ܺ߷=�a�;e�ď��I�B��nތi|sv�ht�Ewb( "�����V	�}Ǿ�6:_9�2���Q�[b�E����g�iC���:�4o-�$lM�T��0A�VxW����Q�H��9��i�>s����"�I���,'N�R������!�&/k��^2�d�D0]����������%�^ �� -��U�?�ѝD������=��i�q2��{�����2�K��;Sv��b��7V���uo���5�im�#~�y!�CO��ٖ���RX��2,-�w���M�뵥�� q
-&Ϸ�,B�a֯��h��;��0�2��ЧŰm���m���c�V�7��ŀm�"�t�+/:]�����^#�9 �"��;0OE��hX�q��)�ڢC�)���s�5������;Hj�)��%k}OIb9��Ǫ���ɦ�E}�Fk$�šRN[�1@[�a��Ԍ��)!�7���f��0TOJ?���	-s)�N�~�ݍ�Y�۫�4�(]��`x؏�L"�-�ٖ��6�!�yXۘ��]#��
>37�1)�,���$��y�<��4?0E>����l!��)h�����O��Љf��=7C��$o���5C?�\4���FU�/@j�~����qf:��(2�T6�ڡ���!��y'Q5�q��2�q3�`��Y�c�����׼�܏1{����/w�"&n-�a.�����A CCU.u�UK�ˉ���6ɮ���d���!¼��r�0z�u\��a� �ܲ�6xd�-:4|
���e�E#K������36h�wU,�i����2/}�;\@��`���L���j�w�~�{�4lg��gexj��� ��V~U^�u�g�i&�׀ӈ�_Xi���:f$�绛�Z>���5m�[�Ҏ���8`�gO�	�][�;�Qg�w!�z��0ͱ�R��H��	M"~�3�	�Ͱ��бmc<:�"�!��S��PQ\�2��/��HA�(�,��8�fv&����(�-���*��X��ٻT��	����3��n�^�9'�`!_wg�g2�c��-�����1�#���V��W9���h����qP�����ܜ��<��2V����t5H0 �@n������y��� C�kr�̒��H�G��.V,'R��$��<�7����Ф�&�0���К������;���7"l)���0�niҹAsOz-淨��4b�(�|�2�l^������}�	�j���p��d����$Oӱ������顃'˓�NF	W6��&�
l^�&�/������q�=�5%����<��3��/ևf=Pjc�e�d��c��I.r���º�_-q�)u	!��H�;o*���h��(��-{��8 ����&/r��#t����0�l�Z���;{)@�.�iQ�0�WD�K/�)�D���g���/'��a�>���$)�K&����8����"��B��頝L��U���I �������_�(���qx�G�&���c�1ѥQ��Y�����~u�����׳�/'-��TS#	*� �o݃J�x'��vZLݾ��'���ࠗ:E���L���lF�Gd����ׂ� ���9�Y.��C�ǹ�ī� )I�Q=��J�Y�Q��� VL`���B3�+�Ny���2	+:����aV���0O�#.�>6"���,���:nT${�w�"��tP�c�s��U�@�:�0�f�u�W���9�_�bLKѴv�9Ug��,2Oc��l�[�����%O{⫿ˡL���9s:�?o6,ϛ�
��ԣX��cD��pv݊p�T#�=�߂�v�T_,��{��hk��Q��i%�F�<)�� a��1j��'��Q��함?�U	��rfj;��I=��B�zs���-��s~݉�T�0�G��M�?G:�U�񫞵C?�W����o}:�yH�%�LK�'-𐛌���,����؋*�/���F1Լ�"兂�V�,�����W.Rx^tT[%�x��nAGNW�����>^�hQӮ,�V�|c��)�h�� t�׵2eڜU�ښ/I��W��r�nLi�!/��yͩ?��sͿ[͜G8��rDl�4�Q���r�����L���,)�׉�T��9� ���39�$�%��e�@9(���&z�p�Ǫ7���,�%��#�Z2����������4aF~p2Y-�M^�~���Tco����a�Id���vx�5���t�j��M�U�]�]�_;2Y���
������D��=Չ-9�m��5g������7��q�/�6g���U��K��2��b!����B�R�ˉ�(+:�W^�f<[O�X�a_����д�d]&h�]?�$
������s�h$3����Uo�oB��aå�m�!��d|�'��خ�������(8��7����ލο������y�M����uLB���]�e�}�H,��ǿ����->�G��fDâ�q ����}oj��ʵ�[�rw��3�*5W����zD��I>�j����ʎ|�{n�T��(]�Y��0��*(�Z�)5l�7�����Z鍠�G� �r�c�{��N$�k���{.�*E2�ӷ$|_n����lH�-&��>F������^�����#;����LT����}#�j��/��m��,�M�`�"c��4�D�B���V�h)��{�(����ռ�)=p�4�Κ�Y��Zf�!qW�L�����1I���q��IXڡ$��e��J@���g����Z�j9�͂V֍�}�e�e�0^�3�
N��*�>z,3�O�ai�!x�1�Mh���ԩ٨e����g�L���d�+3>A�P���v/�8��=�*~":�v?��,���I!@$��($�o��	���h3��_����Ě.�<�|@BQm3t��pǅ�C�xld7U�ݠ3�� �0�!Y�Gͷ`�ϵ�#�g�Tj���`����K+��sQD����!���"��ݢUA`������JY�����n4���#Q�}\����͝��'[ᱣ��,͡�k1�" �i8��h�8�L<� $DC;��c���Q/^+fuH�Y�6���.�B�1p�߆�YC��G]������������-L�K��B=�D�e��s��Ήw��q�s�ά�#$��q��!�Wخ���is~��ٯ63}�&&��~CT'UɪI	�*����_D�KB�
�Fѡ��[$��V|FX���\��]�b ��K��V�S�F����K+������C8����P}����ؼ;��v^�>����KS�%�w������'��t�[�L��Sd=4�آ���i�-LD����6fg
�]6!Y�[���#~��O�ׇUw����s;-1�gBt�y��h����	b�l։Jo�������H��c��3[�]��Ao�Z'@�X����Hrh{R�駂�ڊuJ�/�.���i��h�3/��ʚ���a�#���جQ$��z�M�G��$�(\��n)�u�T�S�/��X��oѠ�b�+h&�.���*5K}ƪ�,M�Ts�@��>��]6��o��C�p���Go���dڭu���~1�,��2I�ۘ�=V�/�܎N:�t��6��i��i�= �qb��&Eq?OkhH���"j���g,���f�~�՚'˕Y ��0��NtKTz�]�3����x���������n�gMD�*i�h��2��7y����Wk:g8x�Yх곖��Uj gURџDXy�N*���i������ʵ���9SF_k��ݵ�_=�w�����A�=��F�[|�.y��\�n��ʚ���{4���K��B���]�h�Э*�XP�{���u�G��1�prU�{(/\
ꟕ��RDK���e�R����_R�d�>�����mP	D���� (����0�b_�	� �j<��4��lF)'�F)}I�<2Yʐ����ь;�H7�$U<�]�/�P뾯��Κ�8�b�k�RB�9�0M��-|0X�=���-�ڝ�
8󤱹�W�����r���?&�+�(��R�L.�+��,�S�P?.~���_�����ş��뻕H�����A��T�����$�$��#���Y�����l@_Vx�炢٫e�S�+÷r�%���9��� :=FO~Y�A�~ykO���E�����g�ȴDZ��cW�ǘ���-��$���ĺ�A��O��̄����U��4<�B�N-�=f���꺏��|�cY�qky��Ұ�4f ���~E�i�)[.�nVX��
ñ��߶ʆz����2S�J���k���7�k����|.9�c�U�7�d�Tǆ��,�Nb0���MK2rڟ,@yrwУ���$q�՝c-v	ɒE���;a�Fn��TPO��4��m��V�\�b��-#��J�3��Dފ�M���R����Wc����@XZ�C(�d	�րK��(������5�1.�#��u�(�E+	�,P����� C� �D��E!�4�)웆mح��L�o|�Y�����6�˽Rx��3�^���QL<O�t���_�Z�=�"��ZuU��B$�,�̓ɪ��^6wca|Fi�6�"�$����3��0�5 j�Og���Q���P���NN�E.�{�߂�ݶ�J�ojĦk

l&?[�X�f�;�V��_�@�c��v��!-��-��9��(LG��Stf�+�Í>Qk{�'�h/W�������g
??�2���`��|�.�o(C�Є�M�	zM�r錍t�2v;������|*7U�8�����9?!�K�a3#۫N��%90	�K�P~�T\�Õ�#��P��{\\�b������-C���_�I^A��Zo3D���>f{P�I�U�?m?Nڂ6�1R���b��F����)��x�`7Iz�JM8HH��@P�����}~�6@�pzY�Ooo̬	%T�	��"�)o`�����6B̓$���[v��+~1�l r�"���N08��E��'ofBr�n�(�<G�/���P�je9���j!]�(�*�3��1����2eU��;�iWH���"�޻މ?���cIYP:��U �e��S�������J��e�2i5��|����~)�e�-h [H��_�Ē���b��kн��#S�:�O�鸀]��(��dE��{��`�	A�T��mp�x�����ߠӼ���hϴ����g�9M�ngn��F��~���L}\R�nfS�QT��S�q���E	�p%�{T3{k��z~�%��+��'�H0c���f�F���}1\	�'����S��73��5�ѷTm�W�f�tP�7�<הd����,��6��k��
��SY"Y�s��K��%��bF�X�u���^�햏��c���`}�O�*���Xk��E���XxJ4��u�� 8����b@*��}�ȼW$7�6����#� �l����Ɯ��cpJ;��aI��kq��=�},�ş��y���RV�a=@8��%��<}�8�ɺ��n�ip�4C2
2���B��(1dw2�M��/u�h|~*�6-&)�����jl�[Z�V�9��\)ƶ��Tud/�(���س�(e���q��m�u՞"���:ˤ���?9.S�A�2����{[d��n����&	�0��I�U�TX�]����\.��)�n5C�d��Au����`�QSAАl�:3?K�6��%|KD>Z�
�M��Q3��^RWk	���]�)��_�6%±���h[�5����͞j�ԓ���P�B�+��P}�E��A�!DN`9��g��}JEP`��4и��3�Rc�`��ȪO=�$I�����S�IQƱ�A���)=��gd�P�D���f{��VX�ZV�xY=�D%��Lˊ,7�G����-q��I����B��L�'�o���bU.�=�k^k���B�2v����{�<�Mg�Z%��W&5��LT�CI> x:�M��S2� T��7w����]Q=4@�� ?����sd�t��b*�B|Y�GT�;Ei��,�FU��ʠ���H�x���/+"uY�<���Jx�K�C`�͕2��[����'�A���Q�@�Ȼ�m�Isg��/b��[0	��0��,�!�Iqğ�Ҫ�:��2q�td>��!�
���>��l�:K��g=��oچO\�=��7���F�����_���An��=�}��|7�X]Ξcŉ��Z@l��'taZԡi�������0tT��;��ZQ����cU������6%��N���J���!����a��3���4�a�I���T��M��{Bo�_h|��vh��E+�!�٭l�S��fԍ�*��I����	o��L��`	]���~z�5٢[�#�1w�$���q��J�-�8P\�P���h��
OzcM�gǦ�F(��u�;���h&�k�)�����4��E��hS�߱����2�%�E*�?I0��S���VV"�++��d+d��M�3�[�BD�r�(	U�:��Zp�����J�?����d����Ղ��v���Y�W вå3=%ݞ�6ķ��6�t�"f�;'��4v0H��dos�!`W*;3j�q���`N�]� ��ƂW
9)����03A������x�x���l6�!P������lr���9��
@�8c����:�ma�^o����5����ŭV���p{�;~MC������I����l�����c\~���YTQ�|\�Ʋl�d�f��!�v��*S ��i�Gt��`H�;�����'�a�(����~ڸ$�,�O���Va�S���; �N4s$��l��QI��,s�L�؟��S��'�]�t��D.��kd���\gnD$2J%�-����TR`@�V��h��E(����l��8j�6�`:�ˍ_z^�}�􅃯���������k����<,C������K��^�cR���ϩ�B�h�����}Q�c2�Eg�(�̌�%Y�_H󌪊�j��q� 7z'��^�|%)�$wf��g/���!4!����<Y���F~V��P������O	x�������U�;�f9X�g$C�p�@�U
f��֏Y�F�˱���r(z�;��HZ�#e���+��ڳn���<��vT��?ި��a+���BP%�� �@``�����q�i]�;�փ�n�\� 6����l��_ba�Q �)fW~�[P�f�l˿�T�f��VoN�k̝j��<�Z�~���jB����!܊�[��Lɽ>�����X�Y�ӄmQ���/.2�-���KC���(��)&5$�����j��"�;����&�ۙ��_�������8OZ�;�81�%�n���!b��+�I$ˍ�_:�隟N���;���*0����P�b�B�((�rwP�N�J'��cߧ��|��fY�}�������3�D�E-�� �)�Mgg��Pun~��|<sC�²�8�h��ٹC~$�#��U�,��v�:�O����m���ve�0��^�\]芼T��љ���@_�o��cp5���M,@���\�7�H���B�)�t�g�(�;�nq¥'׹$���n2L�]32��l�iP�3�PuE���a(����g��5�$D��zKm�wQ�i�o;�Z��l��L���n,0I�WA%m�f!����gJwDt�B��=��|&&�����q�;� �e5v��(:|�B�^����Y@:'Ǡ3��sy]�L���h|�Z�u��v��g^Xl=�r7Mo+����[�νyeq6vu�l�N��a��S�@�;��^Zݞ�^��D�� �O�:Vb�wI�@r�� �x�ސ��p4�x�[��;�n\l��N�fL��-c���$�Ɉ�ko@���|�(����c�N� ��l���ˌ{]�?"��u�#U�o��g��ޡ���j�Ṍ7J���B�쑩>��{�nb��Yr����o�ǻ�F�hX#�~��6�IYk��G�9�LHi�g6 и�6X�e��u�hcc4��U���"AE_�QQ�%�5kp�;�I�aٟ��~�6��Φ�����6��j*��
�ۓA�m��*_l�ƘA��:��l�] V�����?ȓ��� ��ؿ,���v�����
P��E1�.R�@z3����ȏ�{T/xf��3�ɖ�:�?7.%�����{��J�T5l�%���-����0�z�w۫P��S��꙾�:m_K����x4RL�ި���`���i?j	g f������`E(F���!��3�p��O!4��[?���)JJň����z�7���S!~�fJ��2D����٬Ü��\�ZY�~Ib��Ge�"4��&D�]��C�j��b��
��/��+���S�_K���+��~�&~e��P��B!��y2��V�@�� �A�ďG;�.w�j��+Ğ�����t�]�j�w-s��G��8��i���2(��]��ue$:��T��c����ܻ�|Or6ʚ��|!�YMB����P��P{�Ĉ�9�m� �w�Z֐�q� ͍b,�p���t��i+�̓:��IU�yHǪ�x*}:&7)��15U�	��K( ua��£CV�KHn���soG��`:$̱�;Xs�lc�m��#���"	0�G�VFY� |�	%I�@��Z�ݴ����cd>���� ��v�?T��-Oֺ0l�*��ջh)RX�C�ܲ���`�N��m�V��h�.�u�+vHd!��e���1�6?��n����1X@��Y��7�?ܮ��E��>y���!8�3;��Xm��D�1 �91}���j�x�K��G���#1��:��+T=@�S1�:�HN����6��F�	J ��y�m��)}�dZ�9�����������G�Sb��_�"aBn;�3��3鄩W�6)D��T��i鼜(@�6X�rwVƤ �|&A:4�X�V>�C'��V�K7����`�D,��!��6X�
��>@|
/nRݥ��x��K��ؾ�C�6N�P'����04�x6&w;J�g��Wg���׻z���$�SRp2��}%}�#�Od��]��.���rd�������=�Z�{�8��M}����<d�Έ���n�/��>j�W����:b$�2&mD����I·Zߢ�yi�U�Co(�R2��c$�0%\��������L�y�q�$�'��;��!�c��I��X�\:��RNS����C8��n�1�R�F��ah��ң�G�-�k����9B��0�%@�hQ7�j����K�u���nR�3|\1��8`n��w08q{NQ_L;P|���1��=Y}nd�����}p�Z�,Gl�hh nt�k<Sw��ңd��A�j�y��=�m��#���8m�Y�G���5�4Kmx�|tK�[��h����6���O/@�ld�q�W�� ��w|�+��y�.me!��Ԛ�bI��U�Z�0ф�>Z��&� uHN�-���K7���'x�W�CQ�`kt�dH���A��3��X5��͌>zkȊ�s��(P��!�=�E&m�^*��n�vq =�����3'��6t/-M�V2�����p�·�5}g]0���0mT��2�n/�q%�F+�ܨ�%�lR`~�{#
H�[�7zhu������5u𽌬�}H�1�[|fmB�5�ȓu���3�X���9�r�S���+4��~�0l.�'}�mK(���f-N-��s�(��N�P&�bп�2�d��f5���I׬��ۙ�͂A�=`j%9��ҳՈL�C����ڄ��J�WTTH(�F�:]D�z)�"��咻�G��������1[�~+i'��?s�Y��}���s���I�/|��O.�]�GM\0m�0Êt�l�i��I$�V�k����<��A=&6�B�(z� ��DCQT�����g���փ*�P���F�Z�q�穢��/�>��Zd?����Oc�a�yB8�Zcm�.�1ۛ���mR.C�����/����!��[W\�ҠR���:���o�`ƿ#��[>��d�u>��đ����Yf��D 4}��qky+�	lo���k�gC��gV���)O_#='��y��t�6��%��8���C�	�����-�.�x�������¾�!�Y�-%�U�	��D���]$���Y�ع�\-�������i��Q':l&b$�C�mD��rvoͩ\x�܏߆u���ڄ�� r���iJU��}0�u"gǒ�$��e8Η��O'O	,m8]����s����/�#��Ō�E0W��*�����F������4z�o��wa֝�z'a�7۬���fusZ���g����P��)�ÛL��\��[� �&�����!E�{�6�_x���(�����Q\�8�y#6�������:��ȭ����k��Y��E�@W���.�8�ch����\ꦠc�z��& �w��CfTQ�တ���qۚiCJ�;^�
:�#�t����"�הVʒqҵ�Xk�C���,�R�y��I����7jQ��S�f���҄����1��Ύ�NdԌ@E)���HY���$��Nn�!��ՃP�{ 2(ǭ�������al�no��R�@�<�]�)%��G�� ;�O��t���B�dN���ݪ�z��"�v���HxI<^�g�Hp�I⃷��5�-�,�||6��%��䖓�Ϩ{{�u��'2�O�d��?��U�mL~�0J�4�^�5��_��H��y��o� ��N�s���R��0�dw*>vZʾe~��u��g���|w҆�Q��ì+Nt��k��o�B)T�-uD	�ß|�in���j��*��ȗC�7w��^ۯ0B�,k��#n�b�@f6�#�>��?�12?*�ԟ����q̶��'��Z�ƞ�q�W�"��W�;�h�]y�(�&��I�b�� ��Gͪ�e�,@��5�n}��e��n���ba�`��/��b���(�U�=�(��lvw9&(揅g6�_+�00Q �d��t��3%\���u�"Ǒh��J1^�ho��i�a�F�N����Ha��y�FU\��*�����/�e;`��6f�֯A�]ln����t�B@��������ٞ 	9�8�X��,f>�-q�KUڃl�%�((�Ԩ�pQ�_��@-�7�%��ۻ\ng��4,g)x�N����m�5N�#>�<i�W#�Cj֞v���o -Ɓ�JaG���p�o��5��p#�ٍ��o�RP���^�vk�
@.ĦjY�K"����Ff��_x�-�H�f*�������=�k�EI{���i�-�aoU��/٤T��W�;��j�uJ��J����0�),��N�aS'\��5��,���"0������w���c�cpG�j��x�8����<�0�pҢ,.m;Y|z���������`��������d�&�W����)m��S�B�ٷe�J�S(y"qnܣ
�Y���S}M�U"��O0���������k�ѡ}�o*sS�Fv�d�R���֩*Br�m�=�Z'�نV,0�����A�,1���E$n���c7Ch4Ob�Ibq�n�9�4�t��B@�U��c��ygk:�hd�2��I̾1� 7x�������/��TMUP��XK�+<�� t�"���W.�� �x=)��Qa��`L��r}�:Sl��5i�4S��ߢƣt�-�-���I^P"i�0����l��SFY��guFEk����f8(�;c�D/�cJ+�T�¼3�J�"�I|E���M���W94�n�j�!�D�ՈW@��)��m��A}�0��%���B����R�w�d�ke�������5χڕ���1���O��6&�!�]b�/}W�eD���9�={�l�)gF��yZYڜ��������|>�5���0]G�pW|�{��~���Hkl����򶼜֦����b����k�4-Z�2�
8�i������A��褙<�5S4�yD�)���g�����(�_F{�<e m��R���ˆ������	�/����L?��6ߜ�܈R2��7�������;M�2������@#�	t�I8�H`�^yt���M���]L
f���zc����Y9i�$��^�#A�AwߣU�d�ڊ3�`�O*���aଊ��8u���"/n����Î��*l+�H-5�#��9Ý^�H^#F{�g���\*�*n������ˠ�8U���h�'0�S@��|�a�2�>(ek���y	��/�9�iG33�I8RnT��
v�i�1KH�w���ƿ��y�6������5�af`�h��l �oiҟ����5>hRg���p������y0w7�V�0��&��=�y�����F�z����]DxH�jDA�<�T���=�:h��j�b_n|t*GqR_��5�Y��^4�O��uQ������Z���p����>�ѣj��6z7�Z*xӓUi$`j��檓-F���|�,��Ȃ]KcD\�,�� ca��7�Z�Gs$��=酪�%=�X5�f���M}�W�|]���E�i�0����b^���ޜ���>r^�]��N�����e�}&�7������� x�Yq� f�
f;2���v5mI����?�Y�p��Ʀ[�0ȶT	� [�y��q1IO����3h�ト�XX��t��W�סU�s�$~G˧�go��\��,�=Z���,p)|=Q�w���@b_c�/;)E=��d��L^už>�9�j_}!Z�~h�e���KLk?��"��)����g�iUv���|kH��T>W�C���Ioɛa���9&�V��d��uqU}S �,�b�ik���"j'j���0��y���3Ĩ���cS(�+��aO%�~�n����fLQ�I�G���(zD��w��#E��*���5�����uK(Ǣmƍ�)�= �rL�cvo�жߋÝ��:#(E
&�|c2_�$K���s�L,;S�z�,4�M�5�:J%��&���W��	 >G�����:�ĳ�.0΂���u�:��"��2���/+ä�.�>/��FE�9I!�@�TM0RY�סC��>7R^v^0��*����^xM��C���K�義��?~7��;b1P���dt�G�*�0 Vl���>��#�o��B���׳����~�K�j0���03![ԍ:�[.�"��KPb�������
9�/�.X���X�ߺ�*G�E����I9#�n+��j��h',wƮc�r�cs�Cw��ޜ��{���C�-k�u"�;5/|b�I8�|��!pE��h��������鲄e�s�wt!�0�e��)%ֈ��m�cŢ-j��U�)���ix�b���˷C�BH�m�;^H�iF���q��m־7-ģ�f�*p���M�������|ߜ�����F�"���s �K��d��l���pP�ȸ0_�2��R��)�͝���@z�������(�����,g�L�(�2���=��ܭLK��:��g�0Б��@����KK��I��J݀m%���C�=����p�r�Isxնp��j��E0���\#��s��eYa�a}�Eȓw�>^!��U���- ����&�q��YpjU|��Rk>^�zTE��3�S����
|���ĆL][ �e+����ud �˟1�K�%7'Κ��jU"���,�'QC�.s@�`�V��G���`/��(L�~��T�8U��A�x�Z��T��F]P�*[���D�	��h4H$��+��6Ts�!Hz�Z�J �T����,��8q�y�Ű��z���O��_r�\6f�n���V�����LI���D��4�����F���q`!��3�_ը�0�m��T��UXT�d��x�6b����\@E .��WOCfɉ���T�vl䱀I���Gwx576�&G�%ͭ��PW^)��%� u�I
�S��"®�Q���D+�7��H�黐�����>'Q��:&;�3����ۤY��MX��5e	k��7��������NB�+�*����i�&R��۷JYl�
e�Vo1�|����:p�!�.�`�e&���*�wcS�zܽwϼ$��br��?�W��]��ݩ҈;�)�!�	 �g٘�kº
������j����_�]�?�=�B@��"dkR��wR�T��i�����m�y������W���}]�!�����-y�2pj���B�M��һ���Y;��z��ޙ�i~���/R����过�x�VT����}�!'��D���7C����-G<�9|v�/���<������8�<��?�"��p��z:'=m�@v|j�KL+�i��Qzb}"�!�&|�;��I�]�`���`��ڈb?�G�w�ra;�z��cl[�Vm��Z�VOΠ�Ū�
��̂1�Ӻ3�5�P��Oe��Zux��02q�)�X�۾�.��Ŏ��L��״��k��j�e�^{���\��@��?@�K��� *gq���r��L�~N�Xh�x�q�P .��RF�,G&�xn�`����!��|��C�^dg��Y�D̦�A��N��%���E����m��8���p�}b[�fsŷwh�����.�sƇ��1��l'd���'}�%2���Ja00�e�	]�a�&�(��+/WV,�.%���ݳ���G zД��~����l����E d"�PY��Y�D��w��`|��ҽr<���V7��=�<A��4��A�EYW}V�/��p�CXa���8*.��f~�՛;�QmX#��zJLRoo��?�,!XU'.fKL8]p�b�G�lĚ�
AM��`
�#G�z_���%�s�:o����,y�W��t,��$L����	��lc!~�����!��<��p�;�3/�٭��ǶGf,��������F�/�~�Z�Ok��stx�Wq�/�$���g1�p������"�Nt{L�e2��.1*�]m��&��Rs��Lre�g�H���9@D���X�e���MW�.�?T��5W��ՃP�PwȠ���ˍKx!C:�uE7�]�dyIf!�����t�Mي��E(A��;������P�6�K�,�����a9���3�����qA|
� ֲ��f�%%;]d�1�1��ށ�bK��b�j��6�9�-�#mee�w�>�at��tTTAi�Ʀn�}����N�����(�	Z`?��$p�3<zh\d>o�luC������{���)���nǅ�+�5����B�N��T�8�7��������9a�1@{祛)/����5��3�<v��s�k�y>�5�0���7R�JPaZ�jk��ƇI	;q��N)I��N�Yzّc���r&�?��ƭ���W!���@��$���*�4���˖��a|s(��������q�TI���>t��;m�m�eF�W9a�Y�Ũ�D/������k�.��o���cN�X�be:qH��A?ȰQ.aM��p~����S>v¿Zu� ���?�هԿ\͵��DR{V�NG�Y�ʛM��~5L���{8��sGZ8��?0����ٷ5y%y���˝�sU�HG�����l/�[�
����}�16σ_�t�Ki���-�0���-"\��k�i7����7b���D����<64������Q}�����\�	�ѓ��n@$ӻ��.�W�?��a绫!��Y��8�ժ��eP�5OO$cu�@֞u�c��>R�(�%sJ�8��-S7���qw��LO���9a3}�fboo�|!�9��ܐ��
 Q�ms�^�_+��;�2��iԑB�#��:�Ї���Zu��͸V⺨�T��%E���\7x�R
+���		����0bI�1ק���5ƴ�2q=��V����Q��^�t~�1f����0V�q������Q�����M����O��:��Z�CP��$H�P(a}	2fl�e9����6�{�=4#��L��K����k�eX�3Y��Mw`��DG����s7�1ط!c����Q1=R�D_�Dtn�	9p@����	�\�LG�Ὡ'v�P�Ղ<H鮘�O�+���f�3�ǎl֊� (V�@{z������Zb��H��`؉�vR�'��9�����[V��N�6us -�C�$�!���*7O��B-.|�H9~b��?��A���O�8gU��+��a�e�SqV�*��L ��}'�K@w%@x��I%T�2�vi^\��]��U�SXs��Jt��^~G��,�8�5�����w�2'�*{#���oл�,����P���[
w�ǖ8�]s~����Qx>�N e�~��qk c�vCa<�tD(?%�>3:�^2B�HY����h�ޞmĸ ��I�ּM���<k�Tr��c���tW)(Ԛzm��O���/D�*�Ú�ယցq�D�U
����e��ҥ��/+]e�@����#eY���I�92tVl����"���vOG
��j
w����$Rf�������$  [��?�k��=	o���+�1s��i�PNG�;�3�33�n�T&˃_�5s�JB����q�����M�Ɔ��9�ؘ�J�Gn3�g����t>A��x�����`��Fv�A	��(�BR��L���.>���Ρ��e��\��w��˂�y����x�v������<
��k]��{ҳ��!X�${�
i|��%e&I.�~�'�n�L&8�i��)�_gk�!��SY��h������D1}&��Y��*1���	-�}��6I���%�nja����'(B5�xYVe��򌤒	�cԆ�q:�d�&��u�t�KΓa�)����y�޼��+��#������:��D�����?�l�
- ��	��گͣZ�0��U��J�*G�a��w��2I ����x�m�k���1R�*�ɧJ����>�"@P�R1��2�qRʒ4��t��*n�����X��fH��k�#�*����||NvS�x�O�a�l��N|��P��7��E_��(��T� xrkԉTݚ)~�}�Uh�H��b�K8�aV������F�7� L�'���',��G�)<s-�UM=��o Z�vA1��jHP���_64�3��/�����\P�/Nꭠ��(��B3?�ɏ"˷i@�'Rk�Q��;�o� ң�cO�Je�(�<�8�����׬�z�./e�`���}��:n%fG.�^����/�jXm�ߏT+�~���s��S�x�vFn�eW������I����	� ��d�LmL�Lc^\��nLq
��D�y��Wɫ�_Ը9b���9������
}S����9Ν����1'��������^���i$C�$CK�c�(�`9��%r�I�;�ܯ`k�Ήx�6ڬ�s�E��Z����:?��\-b)i;���X���΃����(l[g�NXX�u�+�Ѐ����O�W��������6���2 aq���mAN����=��n#�$�O��*!c���ş��3Σqy�T�R�$�Zu:�����-����UH��OE�>y�`{�W�o)���P���+Ŧ{*�x��-�I��tnbT�F�`���!��Bl��}�0���H�*G{���?���a֧������E����Qh�-&�:�G��ے�?�߹/���=_ZmXk�O_��Vb/���xq��:С�P���*G鱳	@�<Z���p�¸R����`�J����u�OH�r����s�aS��l���X#w�i���ji��x|=b�!0�H����E�uI����EE�w®q*?��I�GA�L�D_�i�=��,9�IƲ�Q�� �t�E�����F�`"�~z�ڡ6�����aT���\�|m��fR\\aՐ[�����1͢��t�� ��pOb�_e%�vkY�QE�q�~sE`�LA�"V����[<��I��R��P&ƒ ����ۗ�
���C���ҰeL��\��z8hOm�F,x�n;s����+Ÿ��z�zeٸC�;�9�!i]~�xMSZ��\�>�Q%�2~B^v���%|o�0L�3�^cM��Z�E�]�r;}~�·���^�Dz��WSg��{�6d�3`h�^�(-�(R�Yb\�ΰ��1�}c���7��l�F�JS�H�͙�$ �d�SA*�b`	���~�>��e�z��cD�:t���aF��n ��L�~��8@ĹKP��Z�|��h�/��\�H�j��$�Ӧhb`&��o0�&>%IZ�;/2X> m������\�D�V-���W����b�|�k���Y[-�p���b��	���?%�fq3V�Ј��cm��ۛ�۪���&��Xs�v���6��E��.�d�%�'�d
Yq�?P�e������F�'���	�#�O%k��nU���o~t��E��E�&~׍��u6T�d0���Fut�����v�mqs��Oș�s���_�����f�eu��:��+,/m����t%���{����O�J�F0/�1��tZ(���^��9�����dU!d��j�~l���0!F��>_�a��R����H�?0��[��O�ԕ*��hUawzDP��3ͺ�
�h�f�ޫ&��k�����b�!�d��T8+���hkO�ӫ0��n���*���#�
���+��:����ж���0!�S���%�V�)�r;�R�K�]ɑ@�R��.���bL�oU�hh}ӻ�"���ub��soC+�����w���ia2�jB
�oӔ5[���Oz�0���î��E���8���|���mk�uw}��=�0z��WF�[�ʀS�9b��(}�#Z�X`��'#VT'�`�-]8w���^��g�X3&��r��E/I�e�4 ���%P_�@�F��[�$� �" ��_6L�u��%�GK2��H3f�)�O���;$��\Fm�q&m�m���$��^��5B,���Ha������ ���f�SpԽ�n��\/�eޱ�-�4Q�,��'�9��j�\u�/���\	��{RFېT����X+��U�f�ߜ3g6�E5�s�{�4}�7�����f�b���wD��X��Mp�4�n��+g��rb�����%C׾U��4)����%�b��*1(�l��s6Ș',JdX��pf�	UӮ�V9*-V=.%'+B���$ʵqտw ��������r1��N��A���EEc�K����K�O��x ib4��%��'�.n.훼 �i��4~;��[j���}�AXD�6J@(d�7��I�Ο�K�Z��>�Yvv"�Ɏd���w�W��r>�Q�Z�(�����}�ǔӑ�&z�����h�}-X�;����f)W`Z2}�)
yѶD������8�!e��.'�3ʗ$�|�1��c�E����f�  �L�d��D�|%�1�Ks�������3�l�t)3�`�D�l�M������sXL,�C��6{�Ց�NG�����1`�y�H_e�H�����_i�0��� ����Os�>��n�.��홅�j�N����@Czx;�7�0v��}�Q�~d�?��*� /�c���+Ίۍ��.��j�<�p�0�L�)a��� z����0kC�7P7s��0�ti@��q��+~p�#𓆂�q��:�u�T��rٱ3$�A��R�tZ�ۍ?(�ųѭ��	:nE}dw�O;ǀM�#]�i��M�
�2i�e���u�+;y.a�<��V�Md����ϔ=�_]GU���1�.�Ԟ��/��{�{��/$HM]�KY2w{˧�/�Ө\o���窓F�'I7x�w���^��܄�3꒡�<ƺ|�}��|VQ����%>���y���-|�m�Z��i���)��#��y�d&��vi��71ݣ�n=�xGV�m�"�e<ʂ<d����i,�˷���H=x挗=�Jw���][j�l3׎Z<h�d�a��I'��<����y����D*#:ԯ�
�j�S��S'j�A�.�4ө5;�Me����moوp�K���z�|���]�^���t�y��.���&��{H 4�M�%��D8}�d�Ћ%�#��n�'��:I��-!�;6~����Y���Ǆ�X�7����O}�����E���u��[��xƪ"$��3���S�Ai�B*+��r*�S�B�F�kK���	
0Z���h$E���zi������}�_7�/R����~�d,����c������:.A�8R)F����d-��^�)�R/3M͍�["�뤉(�Ehr#N�y�RɎz��o|+@���a�(���L)%�ġA)oF�c�k���;�-���I��9o��Q^��t�R�<���U�?v�|w�Wӽ��P_$���/~r߀���\o�iH;j7����DL	��W���D�x��ytP
�f��IϘ��U#���7�W�\��Ru��D��W��mC�
�����P���������77�?#Y䖅!'.V�;6�Sl=�U��]���\M(-�¬.�s?i���E��i!�1kA�@_Od��|dܝKh �K�ry�eT�Y�Am^�Z��Xg�:	��lM�[�z��>�VY}Hh��UbP-�X P�|�'����JX ��K�Q��%��َ�����>��&ȊSP
k��/<y�,'��a��SA�p6'Rng�2�3qS�.�_��ë�Dܘ�����C�+k��$Gxۆ��N�&��WSy���Eu��i���=v�/�����=�=����|s����³�v zl��L�ö�[��\&+pCZȫ�gVX�����W�f;�i�+�;D�,
���J�u&ӮyY�Ĝ�exiM�M\N=>��8�w����I#��촥�w]�"���>�����f\�@�`�ɬ�w
yڈ^x]O#���5�W��f>�P���:����]����*K��}����q$[D�9�Z���������䂁�Z�՛m�B�Lc�T<��>���ԛU���N��|0}�ך������������`V.�������t%� �w���S��ju�:�]5�E��4�j�RI����TF���9�
�M&VM�.��:���R_��]��Z#��s� �s��y��s4��!�/Z���^<ؑ�6�1��S��쿠�}���K�c⣏Q.�\�]"�V����
̓��C8�'����T���#
ʪ.�A�a�4
l��z��]�A~t\X��P���;韜�J ��/�������[�Qe�-�U�ݵ�T�!��M�y�	S W��|�-�Xa�S29l�P��+Y�����*�x���q"̋;������mϹ�I��D}����`J���i�2��j�@*�ˠs�e��䍅�*8�`<�����5����\��w��o��MZ�>���-�l32�w�[����LQʫ��B+ (p��E���D8�Q������)؟���~
.���P��?v�Y�(��:d��z�R~]�]Z�y�^_4~]C}aZ��a'�\2Pʗ
��Ц�~b3wo�c�����H:Z�YX5�v�xܾ�?	��X�u���RXk�M�l��]c��Tww%�;h4��M�d@�φt���<�v��p�05>�%�hŴ
��Q
Hlvȍ�ԉ�'��*�h�L�A����L�����}_�u���@,����:�����u��2�;hE��iʗ�.̗�2䲈���AxM��g�U�+_?峨��}Z����u����/�mҍ�adT��B6(AO3Pu&m9��G�W����%>,	s&�I�ZW*qr�:Al覅��[�M���.H�̀���G4!���!8�N�����9�q�R�ʻ:��I�n�/���� !�1��N�fDe1��J�E=���f@�}�� �񅵂AI蕑���~P��[�a����x�(�>�J�<�B���RX����+��w�ݵ�� �@ߧ�̡c�*hCz 5�X�?��J�(ta�$�7�`�u�@;�(�[�+y�<�o��!�C��tg)��\ӥm�Gqe��u�G�	,�|0�(AB߁�[�mX.a�>`�^?�W2%�e�"�r����*o�0s���{c���Œ�k�s���V�	Ek�7 �*f�˺f��)r�I�8���#�D���V	��^t8]�I f���*7w�p����8/9���d)�+��WvcM���^َ���ѻ�����Z��(�[	M�ފ 6������V�j�<ԭ���uE�� A>l��yT��βZ� ���H�����ꞈ4�h�+C��8dr��F�X���V�T~F]����/�ɇ^���yaԪ$ѐ`"7��>2�&�:Pמ���bV����\mp�]�p��Y3��o�"5�'v�z�x꜐y�$��E0�q�3�y��2�� �|4ks譋4��x�g��(fi(շ�{N4�z�z ���1�RJ�R��{�?ꇬ�q�uaH�Z	�a����^	�5KrS�1�q띅⊔�=:��,�9fY5��&��'��x�p��0�&S[yD��d�K\��*���>�
]�YJ����t�9)�o�P��Z��Y�����mY��� �-ڷt[AiEB��G���9s����l9��\p`Q�K͆Sw�����BBњ�q��W���>��&4=+P�V���hM4�e2�q��.����E���4����Fœr
F�Uũ����)1;)���v��43xvz�h7��F-#�����n$�G
��t��͍zcE�zy��.�f$2Ϭ�S۷﬋u]��*Q�B�� ,�۞&c[���ƳƸ�/�=�Hw�9��^CR�3�����#��t��[���2��&1)sր�+10ˉ&ߏ�a�ᩮe��p2�*v��G�_�x� :aT�b�!�уתb�L|ȁ�tf�X7�m�w<r�y�d�^���&-���ם�Nj�O���s�[f@�����_�ׂ��	8������$n�V�B��g��5q1C��:d��ݓ�B.�p�N�#D+D ��)/]��5�!*�=����x��dN�ՠ���^���Žs^d��:�<�MJ���-��Vm�\�K���Up��b��>G��?@0�4%?����5K���-� �� �k�9[
�X�+2���T��ݕ�-�CT?pw�� T��3{�N:�/�h�67�+��'/R��Y��Hh�&�r���e��!��p$U3�XT�I���|�\D�r���S������E@�`]�&�zoeEX!���b$;�w��+�]���R������Zt@��U���]���:���w������r������.I�StG���g���z���!r9C��ai�� ��@,�0I���Qń�ggΖ�BBG�u���w��c{ǿKϨ��O�/�"���k���`�)���T�ǳ�P3s<z�l�s:>&��e߆��n}����$"R��N����D��P���ّ�� l��8�}r{T�JEB:�H��k�?�0@0��p��b�d�H���\�K!�d(b[��T~n�a�ɻc[�|ۚD�S��3՞P�m���M�2͢`�.qKl9��ԧ��,��r��͐���,Y�-i�s�4 �S��R�g�A�N���k��U��?:�o �i,�1��	�gt��$�7�G�i8�n�=(����\,+�+�R�����E}��/=̟<^<��n�&qI��=WL�)��AL >eQ��zˍF�6�2Wd�ǃY���:[��������g��,H0��tfy�/zc	u��%���˹��G��km�]��ǣ������5� A��G�?I�� �Gχ��r+^��).<h�ً�����2N%<}@NI�kF�;�s��QЪ*��4H�L�ɒ!��b�>4hZ�Ȩ�QȔ.&��y�bݤ�U�:F.�o��L�nD$ [8�7M� ��j��uWⷍ�,� �8�
���b_�B���0����1Qj^H�U�~L/��A�1����ђ���{v�)VCO��r��r��$�hZ�}_�w���ˆ���z����Օc���g�G�Bd4e;�e�U�P�р���@۴��-$�&'5בʈ�^��)��c�w����*=��V���c��H�u�xe�����`f�72*ր~�O����rN�6=m'[�3�:FIP����i�U��݅[�Q��2lb��2�s���ǵd{9�q�i��|]E|�J�Q)�h�sR'�cx��;�&�H��O�J>CP։��A�0��:x�b$����*R�b.Rt�Ųі>�H\�~�Ę�f�\O��v �pͱ$��N$�~������<�~[��8��I��/3��-��Yj��"Yɟ�kX�{�^ц++h��x��'�x�z����&6 h ��j3sQ�ş6���0��	�uj���0��=�Ӫ��Yr�a�ޢ�*��{��N<t��c?�a/�� �{�-�]��@�e7-�ߞ;A���g/pp�~1=ҴO4k��`�\�c݇��xV�Ӂy�	R�2HTVM�st����NB�b���Q�-�}� ߏR�P��������&��_K��s*OA��8��,E�����kgjWUn�Pa�l����sć\�4�"��Ӻjc\G��U4X�ۀ`�ɂ4�y��� "~0��|�j����jӣѴ�z�[�+!)so�v��%�$ow�j�f�.AF�P#b�XZD�1��70�Ƞ�z���J�f��ɷ�4� 9��U��Ȧ�(Μ���x�#m�Q���~�Aŵ(�J]���;Wzsa�?&�����d������i�#X�
�-� Ǉ�O���r�<�	�꛲�,f�?3~yK����w*ui`����0�c�/I�XNKJ/�
��4�C�3믙����{ZD�3B�� �����>ԡj�M�v�x����v������Aє�͐�ol�O^�GBc���.*с_���Tc����2S'��n����]@t�XUI�p��O׼����8Y�2Pb���7dw�~=��sx1���TY�"�n篘�6m���
�p�[�3�rg"G,#�6�S��8�,��*]�������
"O���Մ�r�}�E�ƈ��}����vM�Iw�H<=���t��4�3�$#�6[�&EZ���w����Þ'{
A'J�c~�g[,D���o���h��J��"�F���k�p�0� ��'I}���3**�������,��nB[�\.Yav͚�Ι�Ţ"�PzPk��@�ǜ�^�,p��<(��ns�%�k�:�&{���^�Ϫ3^��[հ�'hl?w�����i��&�u{��! �;�d��h�G���K�5�IF����<-�}�,o�|ke�F}G��ѣ��&�ۢ9���}��u*�������z���.<�/�4b�"�ϐg4�>@J'փ��U `��%k�j��۳����.1dY@���R)�)U��M��E�]��UX˓%��5�F<��C���S�W6�ay�7{�,���ﺳ�4�C"�Æ`5����xn]�2K`�$�x��6* �: ۈ��M��=*n�m���t���䈉��/����b+�����t �����U��N��3�S�
�*�(��Oo�o��M���$�q^�ȉk�)�:��Dߛ���P���bm��|1��������@��V6՜��F��!֯�T�� �t�`T�z^�ZϷ/��1��o��\O���)�(-�0�����m0�2�[bq���3zp�ѹ�e�Z����!�Bn.�9����OT6&���.lavx(��L&��]6����kNΙ��k2�
kj��p�I��w!wdr�� ���"j&�f�_J}7@~/�9��=�׊h�̌���N=Jt}�n"�.������j�@�F��d���ML��!�W�ee�U�yA�kE>����F
��g(�V����#�20c��#>5h;��a�+�|�R{X���H�{'f]0�|�W��j�n�@�`�����Ssp�����V���)���n�`��C��5ljeW3��`�5��j4��Å�����(*�Y#d�����Y 4#Vd�;Yn� v0[�(��넖H���\�US3����I��I����H�:�\�	q��8�	���IK�}�U]<��@�$qy��	�:��z�[�~��0�V���2
~�uEu��A��\eh���yp��۫�`{�T���,�.�b�L���0����a�ɼ{���f��4O3���y�����cB�5?O���g�q��Jơ�+��^��l�����e�tI��X�_���	Y�y���{�~�V@�Wl�,G99��3k|8����ۃ�L���ag��܎ʞYY�47�&�8�^.�x��/E� ����Ȼ#U ��Bз+�)xwSB�>ɨW�fut��$�8�gB���EGB��7����$��¯��#�����2�&'�~K������u�����D��W-�߄����ϣ���\��EOm'��Y�����:�\�C+�a��0c8M$�Ħ[#m�w5b�-��pM�&.�O·ÿ(�f��Xų0jh+��u��=�v�)�E+s��K���3�y�5�n�h�׏8I�����}�=,>D�;�����������a&�dƇD�����x��O���U��D�#Q�=�����ݟ�/E6y:��NɚljʩE��"i~��ۚ��Yb��1ۄl�!��P�Ĳ�'z��Aξ���bg���s�H���D�-1�ĭ���o��;U[V����Js��=7��Q�������	N
�b��G�,<�)��^��x��a�48����r�B�}��k~F���*]��Pؿ���wKc���rx�2�6��S
K�am�b�џX	�6�{�߹��Z�~�'���{SJ/;���k����ԅ�����[���Q=�8��N�Nn�&:/W[����^B�E5��EJ��a��iEJl� ��[;��ID�&x �Tt��I�S��I��g0�$�L�5��H����ɔ�PH\�f��*^�'8�`q��'��tX��C����S5� {}w��/�y�d���b��[ ���#�G/�Y���kx��5�=�Go��X��������
6z�g"�^��8� t�9��PN���p��qε:�z+_*���=�����,h���b��$&�j�%.֭~bp�����6�GU�[G<^�a�'6=����6�Q8m�X�˿=�&�t��Ľm���,�\�̃��Efy1�ykxЉo�1a� �z7<63>b��a/�1��bIA{4ӹ�t�L2*�����b],9����Pl0�jh��K�}�]Uq�>;Q�D������S*E�W��HW�Eڷt�I��f�_�@��z�4��c�
�ݭ������k:@�x�bEz]��\S�� �ڄ!U�A�h��@�KfN�G�[�A�1`�\����/L"����S�I?@����J�oT��r�>��D�9��	~cG&�����0yY��B�p��]�QPLR,�>-a'ř`�;���G���w@[<~�����H��\����Vu�tX��wEW��89 �W�����݃&1+Q	d����QW���r�8���������MT�%��?���W�mI)�o�]ϱ|=zm��f	��� �����aDi��(%�1?�_ޛ�����В�����.ȍMK���%�Z���7�]F]�Z�p����Da� {�_p�7�G�:�oW�w,L7�5����C�	t��W4��`2j��כT;�-�1��k����>�I�
��W���3����mMI,;֭H���#(ѱ�wz^��މ�s W�q��.�K+���j��� ~@��J/C�XzU^�/�[>�EƱqTH_��������Ǯ�����N�!���10����7M,���xG�_^��e��z��1JW>�(��M��u]�\�G�	~� 7�b���2��`��}rV��%�'�6
��H�� �G|g��?�¾�NՇ$����V�q5�C��:���Ϥ�����4��a/���z�H�L��A�˖(�Ъ=m1V�Z�&C���T,9�گ�7ޒj'�mW\쾙a�?Y�\2!i��pD���"]���Z�#�-bU��
7�i5H&	�҃�1��/0|7���T�,J�U�sE�5��˱���Z<���=�T��]�L�e['���j`F�W�՝|��?4�ȗ�K���<�oM�Vǣ;r��ly ������tĒ(�T
�!���h�Bhπ����o#$cR ��^�M��{k0�o[`p��F&`����ϳ_� -�.�<,�dMwOR'%�ִ�s*�X�IC�D���Ԏ�F2�Μ��ք�D�uz]%C��I��h����!���Ee��������gӁ�jNi��W�ے4��Ż_�7�}k��E����gw��Ͽ�x+Z�fb���l+�@s���p�"�u{��r���MM���S�9>�[r9��eV*Ň�Q����/�>�m����>Ar�˪��/�ߥ��2H$>�$�<	%,Z��{b�#mi���(M�%0�Ą���=�L��mqI4�ټ������5m =�������`6����G^��V>��l�Fɇ�)�K#<E�7\�b>x�C)���o"�LYTO���G͢����z�9�I'���@l.(Ξ��v�C�@K\��޵�5�4%^�T� ۹t�lB�孯�͈o"��������V�2*��'0a�N9�p��V���{�H @Fȓ�{��|i��|v�����Sך!��ڧ5�,JG~��T��?��i܃݊t�U`�i�}��S^e"�	RP5I�j=���e�Ν�/[(���)=ڝZ�x��+�w��w��d�����i�ŭBa�T��! 9z.fhŌ$3ԹśҌ��etR����+O_ NN��On�
懢�C�١$#H]u��*�TLN��6~Z%>?��l����8t�>�$��w�>����[��!D f�j��g�ٗO~��z��]VM��Y������TD+����������#k�yb,�ުm�룵���ޡ+I&�;A��Z�c9\kC�����n�Y��iD+�/0�-�$ˆ\Uk�W)_��^���x_fy��V'L��qE"��f1�	p�L���(o[�}��P�OV-�D���;����Z����~�c���?>��l'Pi����`%����Sm��q?�ʒ�V�,=3Z��EV9��T��R'2�@��w�h�qr;�;��O��B��s������K�k�.jU�ş�U���w�:ft4{��N�@��H��AD����Q&��r�F�T�Zwဇٕd	��8t����XbNOF5N �31�;i���������daٚe;�d�0��[�6��|���u;~��>�����P�3��ק�y0S��;��j2v��x��Ȝ��ꓔ�H.� Ir1oM��]�y�f��8H��RЪd9���D1ֳM�
��ו{��e+����W���7NP��N��!K�u�����VoU%�=�[<r�[�u�iQ��C��i1��K(����(s(S�c=$��"0�٨o5�*Z;� �'v�R��R�ׯӼ0>{�P#�31�o;�Lu�f#��.�]�T+6t��L0��n���.d�@�f�~?�c�-�#��Y��
��k6�8Z��������{��f.���c�: ��Jydpw�5�a��5J��]o❱Al���'���ϐ�M�	���*Hv��?��,/I�Q��v��w3_˵��N,���B����D �iyۛ��"\�#�9׆�ƃ��a0��ˎ�>k�й>נ�W���������c�"�SXd&��(
�>��Ȼ�@\��y�[�����twb��h2+_�rA����_$t��r���cUXd�*�����Ic�Fd n���s�cC�u����<�3f�h�(�XR�6��U��D�!��<dA7(o�
�U2�Tp �9~xؘ�!Q��:��/�q����_��������'��5�t5{ǽ|��j�N��ső��씷&��W34I3�),z�`zt�� �p�C���>3T��n���QZ�Χ��W:�ċ��̗[Uyf�?>����@=bZj���2�e??�'v!�:�<EKD��G��WHN��(���DhA��4 ���V�T�/{h~Ш�S�w|�dy�Ng��n�s�o~�(X��&s';��,���}5�Wۢ��OnGn�T��.�f
��sE������ ��,I�8�[��HO1�*�sr��[w��!�΂�@I[�`�JU�{������)�ɯ,2���1��Ur���u@P�[��,��Ap̝U��5�VPR��r���Ӳ�GD�!�	ZHY��a��4�!hld�¬�f�/e���zh Sj����,�¸�����8˴�MY�G�i���2H�'?#,w�J�AQ�L���~� 6�s	�u�{"fI�q `1ҎZK�;��3W��\�4=��y�O�n�c��9��=�'��I��l��=�DH����Hwn��;#_�ps����iem
s\����i�%� �J�kx�#���W�
@�@�lH�"Tn�q����9w@5�7eG7y�`C�=�n6��|%�tZ�d�K*�Ġ'I�u�7~���H$FR��x2l�+�.]�ǂ��y|���M�s�o��5rZ!a<���W\q��vJ�K�)Lz�W���[�E~��D�.�v�PWf�!7��ލ!�pr��}��`����Fm�s���JQי��࿎O$%x�m�x9��p�#`�UV[,_`�'�������Y]/��fP�1�<�Ð��h[흆S���jqJ�)a?�w��#�p��9"~Uv���
��G�:-&,$}����`
G�HWG�u��1~AoT=�]��m�WLm�T�W+�j�LpD<D+�?���wM���$����h��DE�qP����b�)�ڏ���xTu����(	`j����Fzv�W���q��8�Dv��5%��d�"�7f�>�t~�5|�܌����JE�
�������`�"
���E��	\���il#!�a����uZ��;
g���Pl�B�ᨎ}T'����/��z�|��!uq�8L�׊�^?,y�DU:��6�L|Œ�"$IK��
E��qz�X�Y���I�!����H[BY��E�aF��1;F�n��Nm{��X�2��s��#r�&���!���0<�U�2A����Bvk�g���3���p��PH��H5xg��^���H�<�J��ր��A�X����e��YLi�`5������qx�,�g+�}������a���wJ��z4Xo��8L<����Խ[R-Ф�5�v\^�!"��_����̷*�5�.	�BMG���p3�ښ�Q�3��tAQJ)}J8�kҮf;n�Li&��M2���C���
�� ����-hK���]D,mH�G��d�H�1��o^�Z�����k�Xtߎ*���\�b�E
-�ܪ�م��w҈'x�i�F�_�P����äf�å�Q+�iΥ{ebc3>��z���������2�T)��G��U��Z�J[$)�sm�imj����!�l��þ<~��b؈����3K�ف:�<<�9���Po~�3'vv�3�N�!���>��P��&��$������¬�`���)�fZ�K.�l�<κL�&�P`��/}t���m�,ll&U	?�F�ȟ>:o-�O�yH��G� X�m9h��L�(������Cb�E���o�߄+j�1��C�7�0�|L9�5�1FZ�/��A�:�_+�f���O���&Ku������
@�RЖB<�|���I�🁠qA�����y;�/��ٖ��F�b�gߔ;)\���A��5~�AʾmNp� j
!7����/ID
��r�0����L�FJ֡%r�A�����������T�m�#bg��t�4��G ��U`P<��H�Ͼ��c�,��m�ɞ,n�w�vNN�O4���K��-�;�Z���F~�[SJ&��(Z�Hl��;og������҃Fؗ�J����:e�ӭ�R͕l#��#�~����N�ˬ�z��$�h} �Jؤ���� m��b�zAp�=@i{�&ڷ���F>/@J��V
*�b�_ �J;�̴����B����OŖ��џ*��dl����_2z�kхK�EkWt5ʆ�Gv�[�	4��~!��C��0y$�J{��`#Q�-������k��-�a�|Tz�$��>G5�tX���d��pn���k������o(Y��}��L�D���9��]~l������O0I��`�N~�vb����#&�L�����i��J�ܺ_�e�w%���F]�χ�܌̮�6Bw!"���� ����CS_<�!�5�h	G��t��]� d>X;�kch������U ��Hܩ���RfRJ#m0���mf�{^��/i-=@�3B�2��T.��-�X/�
��K��Y�����W����?�%D��9'��>�c	A�a�%����dV�������p#R�!,1��Ȗp�/]5�\����� �1
��ċ8;u��.�9�0�!BMK����4��C��rC_�k1�N,/E;%���I�v����W�5�
��\�
ߞ��N/��}5h.,���։�v/�$�gY/7I�/t<ws��qC��
�E����ʚ�iy����LoWz�~�Y��tW�.e��B$JO9+�`d�F�]��ĐC��~-nK
�k#���3$&E�˿:7E�	��$ŀ�|�YH73��#����Π�.Z� 3a"M���R�P��ψ��HA�a{W�
R�G��9��D�{MH+5� I�������[�<��G�~�;j����S(��'��}ڵ6_��8�#섟=�ap��u�U�Y�R�~%���8s.��������ǒN�P�C��py'�8�s?�[��F~ʺ �'( �}�A�g	p.VI�?+V�|�3 ����ݒ�rgɜ�EZ~6В�[�;H5 I:�:K�yGQ�)���ܒ�w���V��RE��wԸĚ���҇"����e
;�����.�x٨�����yݞ�.j�G~�!Ќ��.o>���Ķ2����mj��e0�A`_�і�.ѧ�?�9443�.1_�8���{�B��L}�Ua�g.�Ic��:'�%�7�M0m?+̗6�Y9�?y�[��%P�H�V���%��FX�����N�GH Ƣ#8�1������	��w��U9V��@W�LC��ft��&�9��V��[_+�v����ȰB9|G�Ⱦw�����=�����j]����(�}v{�{`'I`w9<�i�ؠ3��x<6���?�\���	з���ZR�(.���qv�_�y��`8�
N(�_D*K|u����YD�6�n��r�Ñ���Aka�aR]۹D8�����n���ɀ�ű8��IQ����e���u�f�,8,��Q1�w6���g�9�&�I��5��rcKn��TkIS��Yq�''���j��!���^7�����s���Zv^����cNcГy��y�\O�Ӡi�ߘ�)	2-Ԯ�o]��&Tc��|��M���<��(�9!�-�c,��{�Ly�=<Ҟ�E�=%Wj6��vw�:O<��m���gt��6/�ӁP�ȱ�mZ�9J(�֨�#�U�;���S��w��^�-��HN���Q���}��#�9�E���+	�]��|��a�Q�3G#\��)�4��c�)^�-�#)e]�ֈ^��J��3?�e����6��B��k�0㕀��ΰ|��?���~�����Ԫ��8�+��"������}�:�_l���B��NB-���9Q��,����j_]�|��zʔN��բ�ʑ=8���U3�ϒ>{B��r^_���~T�tUq���bk�L�a��.HaO!������FeIx�D��ɖA�C �ׯ&DK���~��p�Č��d�(
��y)7k�����n��a��1��� ��j�S�6<p&l��b���2��h^J�<51V�+��d���]űT�(����<f�Ċ����z�G�=Jk��>�SÄ�>��`��j
�Ȱ�𷭯ȩ`c0�e�]I�ol���z �ߘ��������<\���uj�^2��@�mJ� Wq�oex���=�.���bO��jb��^n�v���������������І.�]�[��=((&��(>��>��~�`X6�hY��Oa��+����M(�/i�^�KH�!؛L-�+�����!��P7�q����[��b�#]t����t���F��Z�y��
���Z�^�KC2M� Bq��j�6��E�#���*�� ��*���]=�Yek�6&����ʪ���^2���e�[ʄ��Xd������X�c��!�Ȁ}�Ĳ9K��
)12K��~���z���#-��,��!ݻ_і#����k���;=� ���p` �w%[�E$�%����$�څ����Ӿ��	pm�氂��P�a�tхx%ԃ�o����HJ���)n��qD�[m�>}^���ѱ.<Q�[�� ��T)]9�~��|4�Ć��_�G4���1
\��L��k�0�����eϚ0���t��ͽ��}���i���w�14G�v� "
��o	������X`+��h��"|1��ՠ�#�����J&i+q.I4���@�W@�x�7����&0�lƩ�p?k�k�τ��~Ϛ��'�Q�����b�(Υƌ��������RoTA��˪��ط��Rgʦs�sf�nZ�8p1)G���C*Une��;�G#'�y1��#Kp�i� ��lE�mJn�FiB �=�
�|'�%Gsk|o"�F�^���GM�DѨ9��Ì��	������pV��ۋ����'��ݥ�D���O����ZU$˪�rw�}O��|r�-�)вWAU��7��41���:���k�����f�՘���r"�Z>�JmH��K�җ�ZAԑ��؋��_b�Yi�OOH��`��5�#�V�@�i�3��,��$�E?Եv�ϾE9#�y��_1� ���K�仙��3�[V��A�s�s*�]13�Db8�[~����E��5��<�uͅ�^���n����s��u��3'"��<[��͓�t!����`��2C�E�ބt���>Ѷ��r���&�����!�SQ��Dx�����#v���=�����䫣I���7���|[�s�w��4�X�|،Hn�.�!O�;�̾: �w�o��b�eܼb,��:������x���X�ש�o��rE��X"��꿄�b�`�&�|2&�nD����M��4[������%P>��3��s��<����(/EZ�ǥ��ҪE�č�/F�I�n�Dw�;���?O ����r�h�6�\�+�Йf�@�2Y�N4�Y2:�<�B����oI�>Vh���F���/��
���}��b榄�چ�X��T��|��=��p�cQ;��^p� �ƴ���<�E� �oq�E腦߭`f=��5΀pվ��_��"��A&y5�FT}���7.��}���NJ���H<�)�k:��R�b�U^��)��%?��KH��r�5�!T�nk �hW�X
]2��6㈞�#% i�;-As�>v:����j��i�?}EV0���,��b
���Z�wKSg�9F
�o!Pi�q�zh�o���:h���՗1�k�ȅG�U�u���y0���m�����ܽ���ߒ��Q�.19�bq#�~��������ں	+I?��Ÿ��
Z��I ��fB^�\�<t;Yz|t�1�1f����`<��Q���]Ɠc�S\��7�#�I�K�/�G��*�$Yp@X´iv���c��o4���v����o_o<�<%[���1!z�S�z%Ò�ˑj9�����+�#(9�k�
Y
������d	������D�$d�C��y qΦˣ�P/$t��wT/��|T���4?j���s�ۊ{�����Ď�[ 
��R�_r����!"W"@�0Z%���M�O~ځm]�@�xXۢ�
VK�Av�����g@��+rih|5cZ�w�/ �'����o��ڐ~l���}�Z������%Wplgp�$$�71��׸L)m'��s�L�<U6�o�3"Z,T ��(s�a������K	{�	�{�9��Ž����N/7}����5��>�[��N˄|��|N����P.�Wx����J�l�d�dd�����7l ����w�.��]I(¡�ˇi\p��C��&sW�!J?�,85�մ����ڋS�y7?�^y��-��ь���96��y�$@[/�L�<�+l(�(�S{g!�"��d�����������ą|��>����͛/�+���'��5q����@P��f���_��V9?aS� H������"������õ*a���:����.8�˕;�#�a���=�+V�2>��Q�kbG朥�����L5F�;�� �e{����v�0���%0i�#�����ی#N�����P��pg=A��
�z<%�t�䦕�e�e��v}S��}
���4C�C�����!��A�,h�Q�_&���AV0�Jb�O�x��<�R�裻1H��#C���{T��tX�M�ިa�_�8z�	P��s�A�������%�q@�qf����HulZy�~s.��43a����a��y;*m��눒Y%#s�,֑�:!0Dx��Yu��
����	e�bc���y�HpG�FZ/�MI����쩆��X��9�U��*mv���6�8��U���<��Yt�Xl�a�'9UV�l�~bU��H4�e~���yM�a���$ٗ��"Cź5H`���I<=ڠ�������BocW�:�.D�����������՗ ]��*��u�G30A��o�w�݋x���h�����R���]�ظ��X�1`�8(:��t*i�� K�LՏ5j�K�ɫ�:dqe4���R2��+���>G�&�G��,� ��F�����=�;��ʎ��O�8�z�'}�"�6W�G�=Fv�W=c��.+�a�Z�b�x���*�v� �bW��F���J�q�ɂ���A��y����9�ʺ�`�I/���#�����|���`9�=�D
�쵇{���P1�<��eR��C� �St���C�/q���Q�E����;T���x(�v�5�	�z�H�8�B.�Ҷ�f�f�o�� }�Y#t0h�i���nigI�<�V���%=��AY����Nv�;/�m�Xm���%'~��������c��"�c�aY����l(Ġrw�����R�d	K;�JH�R���>L��G�F�j�m�xk,9��Y��HH*���\Q�&��<�tM��)�#îE�E�r^b��9:)�N�)�K�i��� h��ٱs�Տ�è��)^l����m(�-i���Rd�(B�n��.�Ld5M
���<�[��1א��È�8@�auG���P)9X�y&�O�46����jJ�,)��Nj����Ȱ>Oei��q���N��m|�ӼY1io�4�;͇�ZZ@+����M���d�l������´�&/�U��YZ�џ�,�����[��x�
�>g^&��7ȄF�����N��>�� ��:*'/3�Um���6����\4b�:��Rr�+�c|�����1JfOS��d�yILf�ʰ�,)@]�y��CtW�Q��������DK�3d�
&z�*I��a��"@f��,��U�w��SC!nf���0���Z{��4I����,�T�s>���O��;4��-�p ��%�9Ӟ�ʵ�wC����=���އ�is�)�;o;�����Y:�@ֿ};����x�?N�|�g��}��?_,�l��G�v�Q�ܛ�J�xZ+B�G?bD	C�L<�	�Ԍ����E�M���9w��z�-ʰ@ZD>��ޙI7l�n�Q��T\t�a5�d������|�K�،��8W�T�A|WA����y:��o/{2�=@d�҅`��u�P3H�J�����w>���>��/HE1KVX�����K�K9��Y|��:�P�Sك�D��Ւ_���������k�%^,D�����g�KWhM�|骋�p5!PWp��?b��� |��t�7��lpRꡜE��.��n�d7&�t-�zbA���v+��6*@P��r
kqk���כ����I�ȶ�#������
�װ<⃖��(��[�î�/�ڃ#�_�x�"y�{��MӭZ��p(���;������iJW�5�OmLKC!�*PuO8U��~���7�CZ>Ę����UJ��_Lp(�w�wx�v>1�˱ʓ��Ӽդ��oƼ�
�Ik�R_�~8QY`��s.�<WM�1п�d����3�?*���gqgboJD�9�x���椚"cmL;�N��ڒ����p��]��1�����U2��N��6�٧V2�sH�î�H�\¬�7/Z��"�sL4'�hg�y���⪩q���;.����lKgi^����}IS��;#�/_��?$p֮_����V�.��`�	�f���@��)Z�9ځ� �r6�\xE��hl�!�y��P���)ʓ�0��)Uҡ�N hJ�b����Av����:5Ø�����E|Qu��y�E��$���H yۥ�i���g����)��y�/�I����^�N�����Å�r��ydLn�(^@x:e	��!��<��k�ޓ���Я⃦]��8�ܨq��T��Ixuzk�����N#M �. ��BwƯ �4^����ؐ�XYL�0�bEG<А�d
�ߖ}6 �*��LQR���� #5��/�)Y�KVR�VǋC�[�� \�;j����f[�^ʞ<�c�j�YD=���f3���!��.�3�Ң(�Ȯȅ�d�E�i[�0���^B6�ڪ�K&��ǒPj����Tv`�P.��I��S|C`NQ_�6�P��B{������S��gމ����E��X������u_44~�҅�����&9@W6��¼��d��n�^O8 C�4�d����<l���<�=�F���o�11�Y����B /���(�|�P'���FѨ�:I�2��ē���gp8��G��E4�L���8��&?_��Uah%�`zG���m0���[����l�=+�Z��"�ml,�����`��%N�`xؚW��j���Mhr�	X�cÐl �1�p�x�L�#_�Oj�+|��-;(	��3MA���l�J:���SP�j.g�(%܄�c۵�b�2p���� ]�aLh�^k?�[<�4u���m��ҏRu���
�*��O�<����_� v��PȆyq���~F�s��Vܹ�#l�(q��@	�	ԓԗ�[Q[�:zϷ���\޸XzkLj�݀Z�F	t��;0_L#�%m�i�#����#�?I� �W�_�/Z�Q�K�z�b֤��+��կI" �3E���J�a�� ����mP8�j��{Mh�K�k��X� �х��/C#�nԍW_b�źc�e�4�?���Z��:�35�)*u��0,��Dy���ƌ(&�!V�e�iBr2|Ȣ;0��~�=VAؗDwT�fS��5S����RK��;��u���:�5A���7%���<��H�Ô�1�Ozf*��غ���������s��'ޓw����_?��v�#T��(���W`�ڒu���g�A�{��q�`]������^�Ǚ�$5|"N~	ީ�ͻ�VC����|�r ��8,���� ���|�1�}ۦ��۪4Y�ofJ�d l/	��Q.���ٻ�W��*ҹj@GC�y�0�p$��]Z�@�\�6��G-0�
hS!�Bș�d���A;E�0���hF�_�	�;�;��)'Y���U���n-�f�`:��vg�+����t�|H��:��j,G�jL`6w%�*�hIrʆ�0��xS.�5\���x"��5)�4�кGR�v5��O೽G��f�,��W��eS��I��<�D���L3�� ����!Jq�C$I*vp-��/}�?+����l�C�T1�����z�5��v
�gP6.G��H֊�=Ơ�p1nW~H�i!�rh,i�o�C����|�z�S�,pY��A�!:�ץL�0�gW%~(���H���Y|��c?�HԵ�D��]�{�����!���o��;�	`�i�K�Ux��FNվ���[�Mߑ\#�w�]�($Z����đ5"�Mr��9۟��+�1��QP����ނ?,��u�4K�0��������X�D�?P��M]��s�x ��h�m(�Ę�h�@D�B(M]�P9
g�[]�X��O�>��r��nj�Zr9�K�I����9	�,���n<ⵌ�&�NH��鸂k�h�Ӄ�6Lۂ������/�1�(�Kq��Xza�2ǵR���4SL�����������V'��h%�"X�6��&h��%3��Y���b�3
i���ā�W�x����D�,��?�(�eTlt, 0 �8#��
��K�QB�x�>�%��i����%ޚ��o
�T��9.�?�Z��0�}��U��`D�"�HA�2&i�6uR���ab%;��|��5��d0��,U
�|���t'^����m�>7�ք�~>8��t�~Ϳ�v�����3ی��&������G� %�+�H�6��	��H;B�|&�$��Ph��7���4ƚ�%W �l�[T���C�n�6�~�-]'6�3�I�8�Aeښ���ad�ӛ�^H⭝o��tZ��p�d0��*��J?]ދ?�R�� Τ�QKQ,�L�#�l\�)8��@U	���+��z�*D��j���o >b��_-�j�>��(�猡9o�H�q�L��J�ٸ�w��QUtK^��[Q�F�Uus�><DђF/Xc��B)^q�ś
�kQ��T��@����<�<YD
�?����f{���K�W�D�h2k_�x���[ ��L4"7}b�H�~9�9������n~�+�}���I�ؔ� ���y:g�{0���2c�
nY����Y�f�h�#08`�g��uA�7��Gc����d4\�vVm��H�[��z
���X|q�&>B+n�۴,T�#MQ{�R-����9�
ʹ�����ۗ�SrԼ4��O��n}���ay���CΑ�SN�/NX�"�~����j�)���-�f��;i��,����vAvkC���G�;w�٦�g��T׃B�^E_�Sκt��8%���	��X�x]�ƒ�����y^�}��,�~q� �K�!FL�-m766���.�fXJ/`��aG�vl��/g�m��J��+�C�:W�/��	r�6��:�k93\����}� P�t����R)��/y�S�s��눑7�5�[<Ys�&+���^�  Q[^�!-GD/��=���9�^ =��|%=sɫ�'�!ko��!��b���3pEٚ���Is��� H6�������Fb�Qc¹���j#�#O9~��ȖJ�O��p\����|7ӧ�g�f)@ }���\T>��g:��"\�F���l�8% ;^E�<�y��t�S�묽fꃶ�k���\�u�D�h��Z�"S�9��@�����UX��mm�P��Ū� M(�ɿ40�q�*�R���=6���Uu�H k�4a阴B�	��d5!�,�.����h4" B*S�J�kg��+!~ː�,���hЌ����R�Y��.�w��Sb#3�@�^���_0k�l���<���u�8���l�D	��Kwǂ�S�l'�Lcs�-�&�ɍ�>;����X��c���F;a���M|^z�	8���[�MR�[��xf�������ۈob�0��=�-���F�<��v���R�<��m�H��/��Q格��9��3�����K�=�����YBC�2��	
�fd/��!-@�N|l,����s-���O�QD<�ox��*��-T�E5g�f�nrj-�l�u�d�F*��0���El�dV!�����:*Xv���
��1�(!]��#��eo9ǃUGa�}��x.W�X������ 
���#��|1��h8�?��4#�����l��A�?|%��u:��H8�!j:�*<�<m�e������[JH.�[�:%^��) 掾G����^C7�8�g�u�k�9 �ң�zM�!���x�D%$Ű.a�	K
��r&S�#L.g`t=fwZ;��� c���Q���\X[��<�~χ�� �6��4OI�ɩl��#IL}qKh�|��v
M�
��shРd�'�����?�0q�ZK-O(d&��3axa�ٶ��+}�ܠ���d�!d�|��Mޚ��̳�c���8_q;��Kʞ,W��};�(�Pܨ�#�Zr�1�aQ�g^���i;�6��=ɘ�p�L(+ʦVsֳA2�̜�
��o����
�+�z�ZL%���6�J�y֕?�@��-�g1׳�!�D5ŢFW�u�y��إ_Ta��c-3��qi�����bFҏ7n&R&M�҆tÕ�>�:Ď�L���J�\O�I��ԍ�Mw �T�,�)~�j��:RS~�S��Sh�����w7jdSR�d�@��
�f��A1@�!Zm��Y�x��oL�\\`�N{�\&��9��X��i�S�z���E_n�t�R?f�фu�hZ��pͷu�=�C钋&� y�w
�rp�j��4���	#t�t����T��,�9z>E_f
v�v��ݿ�������L;C�k��Q���� �̄�)m�����T�l�b��a[���V�L��Q��H��}d�2��BFv�^�u����y�<���e�-I�gR���Hf�T�uf���n��"	�(ͱ�^\��JP��ԓ+7o���_=��X�OG��qo������dN.�U^�t�/�&�I*��&��_����:�̼;q��7A�ޫ)���	��VJ-&��c�!����:�P�������o����������lX���"Lٚ����.��K��7�8��oiC7�U�h��n��!�\��f���<������.j����`����͆s�0C���EH�F���]��q�����ZP�O�Wg�%����w������ڕ{������G�z�ɺ��-��0����ְ߲^���G2'V��#��Eu>q�;,$ǯ�Տp&�u-LL�_
�^�*f�i~T�xzR0��>��L�H�b�^e�����6}^i9��\&�C����%�Ж.���2hÉ�� a�~�x$����J�H���4��Hn�o���_�?\צD��׋��4W�g5�$(��v���B*�Y�s����~Q������tIx�KC[\� ����!�%�Y%䕘�P��O��$:h^0���E���,f%:D�h�'g��o��閺fC��Z�||>�87�� �[�F:f����h��I�q�Lo� Q�D:����%I����ۮ+��gD�"�Z�����a4i�>KJD�񷍭5�uG�@c�����#E�	Ϋ�hN�ۿJ=Un+1��}N�Ι�o�n��ݕ����"נ�� I���Y�6
mg�2��Q$�	9�/�_�)n:c��ly�	��l���������XV�� ���1+�h����E��f��,����ϐ���D_���K5EvO��-����2x��;/��ܶ�����N@�kvsij�����1_/��1���h{^.�]�ZpdKկY����ϰ���Nw&����#�+��б�����[�Ͳ(�DS��bʱ(��2���/'�i�/A��vvf���=�ī�K���,����{��t����ؒ��^�H%ϘyY�h�\
A���(���`t�w^�������)�K	�9��Y����,Վ�z��*�yf6��]����<��Q�4�-����B�~qo�k�F����2q�Z���^��B�g����iD�Wp"8i�vT�����C�%�X�$��e�,r��	�>g@��)_B�0���I���
ɢ�W�YS�-,q�v���S�GsY���;o�>���@����_+�J^��ת�B��@
x�>��P��9A�6%�{9��d>���1��t$��u^� ��������y)��7�7�$P(�C�mI_����m-��	Z�w^˒���Ks^��ď~:D*���wn�L�T�O�N"Z�=��JW!�d�S�xS��ڧ��${?j��;��pij��v����<�R�����ۼ��N�:�u��d��zםD�d�<T�_��9�+���{���h���wn)�ܴk�۝�����i���TĩVkU<z'ԩ׷�;F����$'ezb&:��"��O�H,������kFN��j��'r>l���������=�YC�.����s�ȯ�����܈h��&�ׯ�g5.�<-�]u`��]X���-�BE[8;FX�㇃b�2=��x�h�ܭJ�j-*�(ԓ�w�(�@k$���X P�H�G�PsSD]��)
Ř�rͯ�dD���:J�B
5�O$�d����Aθ-j+�*.����}�=��P�m&E�7׳����D:��:���(�	G��ao	ZN���S��t�_6&+e�J��k3�?���2�9���j�����b�6/��Y b�8�9_������4�c��x�讝�i���*�b��}�#ļm�Y�hDQ���RX����Nr��Y�D�d����T����*��@���]B�\Fܛfb�x(��;k�f�$�DH�S^�=U�`�SA�(lFb�/,�n0�'�R���a��z[��/��:��;�3�F��Q/�q�(��Q���\N'��Ms`�2tEп�̄�F�Y��8bk��E|�ꁲ�\�~�!2��͵���W|�`�ړ�Y��dŰ�Aں�+�;ӭH�8����Ԉg1��O^�P�����U�����=X���ij���B��)a�$���EY@i`�T������'k��k� 9L��/+�S0�b;Uء�n�:=bv���:������Z��O[Z�A.s���L�~~�t���z��r:f��b���5z�(T���'�9�G�GF:Gm�oWp�xmeǂ�F��^���;+��8YW�� ��4kZͨ߃Xu�Q�E�r3�D�[1������Ք��j�3�����_u�ĵ��C#_�2!�9�0�9Ŧ���/l�G��sω�΍�P�`Us�ɕ�d8i	�1�1[��s��}�㖘���U`���m&��-��4z~�!�[�=�M�����'���*�ǋ�|�I�i������SSW��u���O�1bHx+
��b��:���\��47� ��" ���m'�o��g�Й��+�N��r�j/����d*ŮN��fQgvm�e{	_�": tU��ǔUm�Z!��p�tt.�����W���x�J#Щ���f��"�P ����z��h��HTA���GЙ�*���x,J�U���������v$�5嶜�1nF�}�-��`"�a��IQu�P�PNs@�#Sb'_S�y)��\�����~C�u|��>0]9u+QU�x[��J��+`ͧgo���1�Ɖ4 ��g��ގzX �F0�w%�E�O�͌U��@�s�w;��^���5T[�<#�g�WRHAB��\2�k@6�����b��)��ΗPj�	����%O�^O�G.7�!����Gl��'�u��q�h��<�d ��	%.�C,���>�D�G�\H������ƅ%��bL�x�w))|���f����|^>f=m��g �����}w�T���wD��`�Ķ�J~#�Ɇ��T{�;��ɴ}�O�p��1�`�$�*6�����eU�6i�Lv"NQ�'����ɑ���I8���PQ�'��D���ʙ���wf��X)}����r���]�X���\�%� `Q���K]�L|t���E=MeB�`V
��`�]�~���O�'����Wh���f�Vݭ�aL&��-�݊"1eM�Ψ}]��Xo�;0bu�O�,�S�ڛ�L �j[q��W�|�͟h�s#�/��.�(�.֪	��J�ſ���/2�&��F:/2��l�,.d�����Sטn����9��)O ��k%��;���R,�X�����3�[Ƥjی����L<T�$���VTh{%�#op�o�	�-p�+��j����DB��7W� ����q��O$U�F��|feLջ	����ش�+�?�\]�Ze�Ӕ���^�w�ƨ�tk{b���yt��B�H�x肻�����=(����rk�&�9��#ѥ����Pj	=�Q0�6�o͏g}��I���
52��'���e4u�-O�ErTŒ�A�]��H;��r�����#sU%N��Μ���!���PT{.3�<���jU�k�4�J��%./��J�c����o�u�ag��AP})��W8�������q0����!��2��`�v�R��懐���z�xV�M�G�S>h[�iS�+�����~��4D�l���2q�7�����R�4r,y��W�v�ɶdvz�e/�KRj�I众�Ր{f�z2�Co��O҆$P�1
k��a�O�:���T�a��LwV���a�˛�q�^� v�?���Z�u�̈������������292f�ƇP��6���.S�B�@}S+����Zf{�	��S/:ւPq#y�<)}��.����h���pV�%y3���W,�J�/�	�,��I�C���26[j{h���21�2����P�y�L��1�,�g\�8���m� )Tk�#�={ �p�k�i.=^�M��q���n�	=�&�&?���G©\��BM�����+t؈yS��>���s�\6\��*���I���^ߣo>,��$}%v��̓P���2�����Ɨ��lq纙�s^28������¨�[f�Y>���pJ ���Z39}X���+�p%:Z|q��P��$NNѥ���d�NW�?���Dz0�f[���+���o�Sn��������2��;���_���3Н=��?��[�;C)?�[w�l���ߴH�U�Y���B+��Ҥ�IB	��᠉�2M�*$�o>�:�̼7�ݰ`��ǣ�Gv��/kwO�l��Krz�SI�t�m�������|"��(un�S��2t�a
����7�FF�=D3�2��I�;/e��Xw�jޭ�X.��*W{����R�Cٺ�ߎ�,qY_-�Tj�c��ڼ����������h+H�`���Bp!�Dez�:B��h;n	���~9p�NN�������/���U�%A�f���k��Ӱ���yryb~�Tti�ܺrc���Z�Hg%�	l��Dcױ��)��OIO� 8C��Cw%7c��У/��0�	0ϰ���(#��x;����J������I�Z�;�񦕠�4'�k(��ھ�]�������c8gnْ��\_e 0|=������mn�Kc����hȩ;���LP+�H�@�[����]	�����gq�w�[�,����l1zT6�԰��'�/�Pe�n7`�Ey����\����v�
{�?�k��9<�C�A>.��l\�5s%ֹ���`�D��ZԄ�\����h����4Y1��Ym��?�4j�2S%V��(�B���������6p� �j�X�^�X��F׹�V��M�17	D��]TV�lG�����]_��?['�O�p'�6���X�M�T�*�h�ԑ-oc�H+��3�2W¸Y�N7[���B\ojH�bK�1�*���\�A��}^94�-�����쌴@�g*�ӟ�����l;ή*/�:u�����Q2��|jJ+����ׄ��Ha���J�uƝ����L���%y����>�������t���8�z(���zW޿'<p>p�hO��E��(m�6�ʲx������L$м���m饖���;��y>���͈���%��k%�טj���JdIۜ�	D�Puk�b)и�R]�W�6�zr���b?2k�40cK�z�$oZ����KG�x�\��3|�@!;����cY�Ĕ����G84�3�d����D ���t��((�.ǥ�B����G+�p���j8^�Ny�h[��%��a�g��b��݋Pԟ'0���3��|�l>>����6��m�_Lp�5�u�B5e���	���[�s<�j�@N��w�xb))��WF�6�h�@G@�63;t�L{�g�����,X��þs���`�G�P	Tv^i�y|S��6{O�2��9�%u����N�9�ך<O�N�$�H�:�9^���7��JΕh��X�-���蹋�c�1��u#����@��A�`X�ʊ�pmb��l9�T�;uU����ӷ1�[f���!��v��t����CU�o���qƍ������c��nHӝR����S�u�1��^϶�V"6���p'���4uo����WV@V�8�KI����9F��֋Tyn�m�o�U�|3�G<��Q�!�v�M2��?�u�y*�yB9�M�t(7_q�9�2�ib.5�a5㮞�=��+�]�mY��Ba46P+`M���hl����^�z�h���^���L��D	�ȂL5�\�m�99T9F�N�~j��_�t���_��LI�S��X��]�g��pn�̾{q�9)��/p'B���2��X��f��OI��~*Q�Ge��;�[ȷ��9l��)ظ��2j?�*�'�	lB�1���
oz��hx�\`.~n�ה����a?�~��YV���+*�_�����x+͋y��4�+���81���
�2F1����v[��!CK�iw�	�6,[:KCxs�MTy�������N���ŦGN�jiY&?k� �/8�U��G��n�T���-����A�X�< IN�/�P���d���3*����C�_7u\&3Q�p`:A���f �e�8�!D�Z�[�~|�I�R��{a%�?� ��?����C����� ?�$�\C�C/UmN� ��\޹��t�?����@$#�׶PpD�E����c ��U�	��0,|5v��M�wf�?����ۃh�%�ac�td�|�b�.�}�J��r,��Tْt�^߇:��_ఝ4d�)�����t�j�6�ܙ��0�X�I׿A〼/+EJ��9��B��S)��1�X���2+s����0d)��Ĺ�7}E`:&�!C��36���P$h$���0ɧ�Wq�W��Gb&�qv����Ƌʔ�K�����Ͱ};���Ѷ9cz�� 7q%y-A鶞>�<aD��?�N�i�$��e�ВE������U��od9�v���֗S_(|oBƫ�����|�a�|��	�d�y����26|�2c���������\y��5����L^��l�w��l;�|8�S����^�7� 9���x2ۆU���Nc: � �!i'�\6��d�5^Զ,*N)�ʻx�z��������P�-�:��������t"z��j�&��}@��eߧ���~9C'�R�
#�(����̎�s��q-��#����:��ǰ�`�	�Y����Fs�&��33*VM���������M��W����������Ȅ�16h�m��"Ǭ[Z*/@�F�1�0�^ᗣ� ���e��Qm�T��U���0L=���B6�tu>Y0�Ϲж*�=��"K֢�^$���H�g�:��G�txs�-oQ�%��o���ɵն��;_��8т�PL�߳��5)5*���4�Y��n��1b�.&8��IA���G�|�IK}�\�" ��rx�yN-�i+
����#/#�^���	����F� �p�ŗ�)��4XP���h���ބ���d���?������?I<���y���c�B�h@b���9��P���0K*���bI@�����/�)y#h	])d�n/B$oГPy�fŵ���o��_�=p�c~����E>-F��x��O�%�D/� �_q�?�F�ݬB�|���*),\�����2��[�iN�g��1�nf8LE2r#�uإQW
��~�B��c������˄]���k���O	��*��&J}�tVx�O&�
��̈́�d�/��d��'�����,� ���ئ^?�\գ���,L0�� s���ي��g�Co~�O���v��S�"l�[Up�9�.��<�����}��ݸ�C��G}ô�x-�~)բ�O[�*8���2���e�4`�v�+� �g�gM�1}�.[kv�d$m��|����&%s�: �B8�8NiP+��W7_}QNf,ьE֍�29��D97k����H]$�I1��^��>�Y��dcp�y�Ss���`�PT��k�.��9[8V�R�>:���;�Xk�e�=5ћ0J��2�>)����{��1���~��Ƣ�3y�/ �˿&�t����m�G	�u��3�r�����Ӛܣ��p<C�]��5g������m�O���#ղ4ݮD���ِ����O5��-�rA�����, ��Gח��r��;��Gp�q;�/�9��$���A$��e"#��}?KL"e�^2�����H�d�{�#D�ed?#�$vC�/��JZ1dS忉�]�w3y�C���B|�����Z�d���^��}݋�Jtt�n���[.��D/*�q{	�o-�J4�s�<VL��0rr�XJjLt��O���?�z��K7�YNڋ�6)�Jr�) Ŭ��-NH3��^{�/��O}H �3����>8ܮ��@R�}2 u�.���کsEmi�̗Tx������3&�׿���W<�ܭC��N,WM�c��ċ�'a�O�͢0�!h������� X6}� �?�K�)��<��y�d߰�kV�_���En��;z�j��&��p�	310<����i'�ئ����B��e�sz $��������5�`��-1v��*[J�[4�S��Q.�Tɧ_�S�e�SS���z�Ev~N�[�àe{��;&H��@yu�*�S���7�ǶHZ-�,�𡽄�5؅�'��0Ix�4��^�;��ĕ�Si$�`��i�fP��QJ���t��4F�����f��.Rٜ9�u�ߑB"to��š�2�6�����"nЬ7���5$T���e�,Y)><���z��g�~�T��b��|�gF��==��#�����\|3��}���b*"���+��5�I	F�����"�Q4Is�����c�0��r0 �SBM>������h���d��V�Z��PV�)���{y���r���
LRV��g�j[C+���mQN�D��1=�L2X�20mx4��	�_az'kV��bX��_jg�Z�R�pa0��-��ҕ�����k#l�L2@a���6�z�^Ƶ��������
E�RD6���vL��e�	Ǿ��-��ǿ�_' ��?H
A���Ht�,[��f�3@`��r_����jmV����bxf����|�<�+D���RQFmc���yK<@´�	�E�gh'�'*Ҍڕ(8�vb���SꙎ1C�6
	G@Z�@KS���}؄�m�5E�0���U���8mU����/� �bn�v%�ؗ%��G���{gD�G�80�M2W��,*�s\�t ��i�Ȇ�rɪi�<Jzi#V|l�X�?g�5.�skt�����1u�<-	c:�����F�e��N3��z�h��5_���K�����&8�7�7�m�sX�1<�z���_Q x��0p���u�bk�$�v�{�@�ᾤ��$�Z��S�A�5<(�T�6�^A'D>a!�)˭�K?b�����<�V_����B�Tx��D5�������OA��C|ZT��e4�V�8̳�a/�f����Y6Ag�p����؈8¿V��O�Ձ�0�;��W��:2��S�$�]!������4��~��^�m%�p���y1oa��rm�%+U{5�WX�8[�Hp	����:Ã�<����˟�%A�y��Ė���b���b��e�V立S�����dF��I����i��Z.)�	�k��9��t�%�'�ӺtԔ�_a������m���!�dUӼ��O���A{��Ϻ���ld�@��P��L�Z֝��'5[����$1q������U���%Ւ�-�i��I$/rАrR�g��̽N�E?�L#&&���B:	�<��Cs*�R� ���=��V��+�0]����c=�bY�>���R/,�F���&`���,$�W� 1�O�doyj̥Ɏ��@�(R9hѭ�%^�0Ι�s<x�
�e5���v#��Ǖά�������!�Q����vs.��ZHY�w��G��h[���������]F�=c���?���T�O�8D}R���3c�Փ�b*�}�����w�p!)��
A���c*�6���1*HLA�a7����6�TӖ�uPD���Mۄ�KP{+�a�;�S^�ew�B��y9�`��*�]up�꒮p���1��N�I�i��*ԏ:JUH�ݒ��"0s.��(�Or��.2Or�>��c��_�^�(����6�,�=�3;�,<��f��E�g���)`&������HQ�q0Ă/N��&�T�i�H�\-� ���f(ڱ��i@s3����c3������o��!��ajR�h��V���Н�y^�����]���Z��-c'�a�?������ܺ3����B��X��A���`��]�� n){M���}䲟 o7Q?i	e�m@��)�IS��W%�FQ웓n+�0���6�2
!�z@�\7���D�\�f�\V��giS"Ry$#�H�߿f9�~�dN�P)�MR	x�{D~RD�<r�{�%*3�SƲ�T�Np5[��5�L%�i:�SB�;W��2D�df���	^sq_4MY��;"3m�[RTq@Z'�5�D�uz���XWZ(/�-����*G�<�x���[n{gB�Qo��ZsM�ai�W�Y��F�:��#�,�R����A�.���%Y7�S�c���ڞ��3=��|�"-���wCI)����������X��שn�U���CA�)�/i��`C9�a�Ua/eȔ�-rfHiSzq��H�5�#�4�#�$]I��w췹�	�A��KC�񦼤�����\���s�f��e��6��.��GS��)�" ՝���p�b^Eq����x��i;'��"P	�'��(�؅�R����i$�w������r�2{�����˫Ǆ�*�g$��H����Y�5�_�r_���N�����r�eR��G*��M�Լ��+R}B�)�a�e`���lL���D�n�����A���Nmi��X�i�ox�g�u0��̱��9�Vwf��[�x�� -��Ӝ2��rG�&�i�!�,Q�"�"�Ѭ�6A�DL����D�����i��g&dL0rVxű��zu�`�n|��b� �� .�����%P*����eLE �n����e�Eŀ��\<QK��P/���7�I�Ca��Lϩ�vx���$��FE���ᒍ>0�$?0#(����qn��$��V�	9��h��I؏�f�:���a�N���U����e�+Ov���-{�d���f� �n��"k�x~���Ϧ��04��3�s�����XZ���ak},�_�y��G��2�̭%�QD��� ܍�Ӏ��
�9v��Zic� �;���eq�ր�Ipy��D]7�� m��{��X���!��sx%}�G'�c��)�!q00ZL���C4�(�*}a9)TǛ��ᾄF�p��A��s�%2��
�
ڇQZ(��nt.lƃ�D6s���!�@Jhf>g�[��AHY?;� o���f4����TF�b�5�m�X���=/ ��39Ώ�� MPc�hTT��Na3��YG��ِjR���'?��h_�Iت�IZ6L|�`�{�V6ҥ?P�;5�T$��T:ˢ�+(�l�M�O�@XV
���|��4	M#j5��pH@i ���Mˏ�T+16�R�Hc�M�Y��%�	>W��
^�2���]�M���1��$�;�@[��tC��i�I!v���M��ū|�V�����b����Tr�W�U��S��]��\�..�A�Y��k���M
��AraY�2�D��e>����(�a����q_���_at (��u]�xҮnK����2���.t�`уT/���f��)�9�-(�ǋ����o��]�"������x�oL�/����rs�T\�.�#��\B�Kjo�fX���b�	�A�|�AOɵW�ϐ�ߛ��a�N���JZwثj[l��A� 4�����a��j���^
��.�	w���G+�����-<jݍX�t*-�Gϼ�A�4Ա�.Ǉ�)���t!�򽃎�AװF=��ű�N�&{ ��y�	c��VH#�\h���u�$�Z��%�<�rv��V�@�ƠQ8�s���<<�z��Q]?���T;+�,}�v�}�*����R5\��#���*1|g%:�w��X�Wx�`�3bøT��6L7*a�{��n�^/����TX˴��V�B�����x�ƒC�%�G���XL ���h�D�w��"A�6|a6���d��J�=������)Y3?��Q!|V��K˶m��_>/!���\����^ʦ`*��cdL�Ǣ��f��^Ө����H�'��y��K��9󤣍�n�������8�C����GBSz1Y,7�|kK��"��x�����50��ۢ�>YE����&�C ��3JSw��vn���k\^/qSd�kWD���nk1�z�%Q�߀rK%Y������o�-1���ǖM��ػm@�y�l5,���I��_�S��Y�ض)GѰ)��w�*�O̵/
VhW�}f�?U���W�%���=zMK"r4�e/�~�Q�����)'�c_�R6�~�;��t�+�Ҹ�n�u��>֪u�J�����5 jKV_n
�������E�8�ɼ��q?b��'b�Ź�ݴf��1XQ�D�zC7����9x���l�*<][#�IL顣��$�Z�R��l�U/�Y(�͈��)��TvMl@M:�'�����{��H.:S�BA�8h&
��1�U,��;/σ�cϣ���c�tmm���u��o�Z����D�`ǉp�M���6�����W]B k�~�0��FO��� �S�=��]�C����Q�z*(�M��a�<ʀ)����n�O� �� CT�~A�`�]qX�;C���+��%=�gkb�	�ۘ,��`4垫D��i�r�g�'�3I�@Pvbt\�QbFz
P_A�e���?tX�� ���϶Q��Pѫ#��{0>�n������Ɂ�$L��j��Rȝm�����>){}&���{N���B�
��ܪ��[����wЪB�L�yF1bTp����ՔQd���O�Q!�K&Ń(���%�wz�g7+�ǰ�3O�̤R$��&��8�#>�p��2`uG���GM[̣Lk ?L�K��	O�5F�〉�:��W5�������5���C $7��v������wqB<�{�"g� �?�ש�>�	���!��*����1�Q���R�)��42���״� �@����g��;a�s;�'�k$�ԯ�O��:��C ��� !,���R�޲��y}�q������,��S�-�|���:��X�.�;��	:�U+���,��BJ���9h�P�UO�A��V\ ;�ܽ�X�-*�e�Oۺ�S���P�.����e[R����ͽ�`�+����8��&}|-w���N\��fa8%~���-z�-��ǂ�h�:8K����/d)� �a�=�x�����hAJS�ؾ2��WV�`ׁ̥����;�O��4O�¨p%t�5sV�tS����L�ˣK@s?��4YY�"���l�Xs"�3{x	*�{ї�-��q�Nu�������Ɏ��9p��?9ɭ@"^���K�d����!��N�-Ҹ*���4&8D-3�J*g�/+%֠���=ͯ䄒���X�~Um���2^Q�H���O�P���O:�E�Pde2�3�}i���|:I]4	�=�)��M=b/������G'��ͅT�╮!t�Ȋa��,mb���#|p�`D�n��{{�*��N_Y�����*��$�8��pL�최���j�W��o��������7?.��vZ~Q,P��'�K�T��B'�;s���9����i@���N���MA
}�	���diQ��)���,�/�UMI�:��_������~q����6H�w�	�
�Ĳ�B�����|q�pw7@J!��^�:�rD��`pq=S�����̺Ou��x���щ���P��d;J��aE�ރ��f8���^ 4��ۛ]��v����=�W���Q	��]߸�u��O����ƒ
G�N'���q0҄\�%�ߘ�2=��O����@3��(>h㾘����l&����|�|%@A���-C\mg\�D����6����$j�%���i�4s:?�w�8>a�a`Ź~�-R��bb��>F/ͣ�%3�3瓑���� �
=T�:0k*�W�5"ġ�=��f�7�u>�[���؍.�d���t�3c׮c�0+uW�'͊�N�س����W�l�Y��^�����U���z����ڐ����� <L����<QOy��Z�Q�P�i��p�c�_[	>�ͷ6�4e��&�>Ǩ�\��E4a�a�gŨ����ͩhK���3S+�&�<�9aJ��h�mL`+zeE��n���6Q�kF�)��{�z4W��i��Ļ�^J ������.��"��]�B���ܧ0�Z�L|����i��]{j������ܚ�}��?���=)Ice��¨��}�7[]�rjS��W��ZDoj�-���1�b��H�vt��&#,�"X��q0�Yt��7*�2v ��d휥�ne���$tc!B��p�k���\3K���0�D�o���z���RW�':9�{����@����`ݛ>I��e�,5�_�O��֪y�d��n�JWB�h.���G����T�S)���pߕ��`9m�cȷ�4,�v�_w�lh֤c��I�wj�GD���^E��ɻ����8���C��#�4�O�H\!�%b��������}�����)��x�@Ҋ�OV��Ě�x/��=F��-5�ll�}������g�+z�נ�k��U_n�+ֿ�Q�MC/�#Sv����"B������J^b�Kb�򉋷��iG�>W�c�Sd���R6��**a�}����,v�T=P)I�U��e9s���=�!�U�7De�2U\c#�
�P΄72@������X�����J��N�����xΫ3�'�E�U��K��O�ZG� ��y 0&J�|  n�c&u����TƩ��jz�CdMH@p���p�OZ����:��.�Ц�t��s�g��4�-4�tb��#@�PF-��t��%���DN�A��|($fqQx�����v���cl�L�b�N��_��~�����U"e_!6��h�<=�[�և�����	"u�5� ��]wn/�:W錄ϓ��������'�J�M�o�cxO�\�"�������}ҙ?]n�Xo֜�*h��&�]�8���.y��e�@�����!�#�P��i�S�4� \��}����������K��	�j	�����0ľ�Xd��d:��\�0~�)��b�T�5�~�Ć�~um"|��c
^?3ư�K��{��?G$$�!Ci�d�}q�#����k�h*�v���P��"�7�h�(�O�{��b���b�ҽJ'5Ȧ��L4Τ��":��h7g){�������p��lZ7W��az��s�i��~X�j�t	�76��el�����>��#*LH�O���«�G;�x�Ƶy�(��&��[_��o���� ���?���ZF�.�Z��&����ct�c�T��N�p}����mV�s��<�%��w	����WB��
#�ѓJ���d.�F�oo̮�j3���U쿛Ov���Sp-�MU�Ϊ(��p"̰aaɱx�-��G��4�e�}�R�ܤ�X�p��v>����xgz՞	j,�*7��Q�C��g��f�Zv�-<�Jp_r=��D��g��w/���:�1Ytc�����8���l�S��2\�M���W�^��<����\��Y?���n�%3��d3U&��n^!�S�%����M���}�`%{H�p�O�����cԽTa�w�D����FAPĄio��&�����ў���}������W.�Z(�&#�⸂�x��>�UYm�������T
��g���u�o�m�\��L-�&���z(��I.?ޓ�x���f,�Z����d{����91׮V;��t��@rPj�:G2Z��Ok�Au?�aU��e4��F�|�wu�-��J�W5LxN��|���4[L9��l]&�L��x�ϵj��~Q��?��}k(1ʌ�������4��%���
��נB����Ml��\~������jiK�M�>~5y��C_{�8Z�qVi��
�'�=I�BP �ܶF��t:;Bx�R)!$��Pg�!H6���"�A��G�m��Vvtk�F6q7Op��e���F,fo�"�D�0z��#����f�VrA���P2����5HL��?�A�M������W��ȍ0���7�ѴO��D��!���S;�,o�W�!\��0�Y�*���t�Gѓ�I��ՏȐY����,�w{�A�E@dJ�]��r�	���x~��p�>��F4�6Р;г��E-�0�*W��i�_=��q�:0ʪ��#���@��6Q�`AQށg^�$����{�ge��u;��yqnG>O�m��Id:�:WV�b\+��$�7���;�ɽ:��@%��ntp��:(V��Q�0-���;*�Jۿ�� k���!��4�2۫鱌hL8������S�f����.1wVJk��ꐧmq�0��D<�<��lJ���➋�m�2ʱ˪�,�m0.˘�?Uj�hp	
M"E�H��"v�W����0�7
��?<h<���V|9J�!�FW. ]��[��}O�����U�#�	�!��yo��:��3x4{'4�w�����h" �?�-x�R�����nRLRv�+�K`M쉐dI�zZ�֔��T�7W~j?�E��.�a�}O�T�����	� 9��2/;/� �cN۵���{-�wB�fR=�C�Ci7E����4(a� �zm1���@M~
��֐]b�K�?xWux_�^0�4�z'�Ic�����[.�b�$���KUʣ(iƏ�u�-DGF?OWs89*5�Եd����[7`8�5{<�&�$�/{��L�7�~-D0|$��S6?�뗕�u<�����;�Q���5�tC4��˵HI�Bǩ�ˮ�3���/"e�)3�2/���f�^Ը@��I�s��g���l⏸�-�J��p�3�>rO��bW�
��a0�P#��3�nzE���{u�Mj}S8�D|iY��C�א�~2�O�=g��U)N�o�{>̏V��3��B�K�����f̼H���ZG�@��bX��S�cw�/���vz�:����1�_�)���B,��
��O��4�T��ͶӮ���y<�S���djx�Yku�Ƶ��H��I�V�FQ�r��$�$榀�ɥ��u�%u��@~��@x�p`췝J�:m��Ξ���uw����h�{��^��LB����.��]lQW�2�����;�)�h�Q�L3%#H"��� �t�	zT�erJ1�z�32�u��<)��G�!�Uuc����_�T�HS<MZs�d�����N��:�A�2@H���,x��l���V �-i��$îH~]$e��Πゔ��5��\����7V^I1�e����'�Q*��8����|�zSnԵ��}���Pv�ˉ����W��:W݉�E��[�\���Y���]�)!��K�"��9���CSx%�\���V��Ť>�5-��X:U�����I
�����0);*��c��3�i�!����Xk�D ^ q��j�ʎ��n��wXvу��;�#��y샸 J������O"����|�r���\,�s&�j�}��C��y������J.f�$�+略D�S�w}���je�9$ �dh�8`��q��֜�>���]BЯ��G�|ޤ5��BgV�����kBZ� �������	�1!fuT'q���E
�6��q!=��-������Q�r�q|�SP�m�a<:���Y]�:}�,e4� E�	OַR��NU��v�H{�z��"Uk�w�] ��HXÐ��)��tY#����o: b"J�xRq �n����G
_pN��ӳ�׶��ڳ�܁[�dB��'�+�����߅�����>��R1�����Kx��֟q1�')��{O0P@��K�.�_��0��+Mw6�D�QR�uya���0��]�]���7�o�6��w�<nH�EEһ?�UٹZ��^k�UX�w|>�Q�#C��e��|' bt���"�����9u85��ml����QO#"�&'��:)ԁP拹���H�ࠣ�k7�+{��b�TЊ�9��R���%n8�npL6`�:�>c0!A_�;"{�jD�&���T�(��fLFԵKS@�=m�d�a�����X�g���*[7���0I����cRU[�g|�{ /�2�҈ʽ���1#F�7e�9:��{��~�V���)	=�a&w��o�}@VҶQ'�%��Z{�r=�v̘\�g�yh8�����
WM�.h )\����ŒGS�J?�`x�5�ox��������B���̾d�(���xt�By��9�ȂM�Z-�e{n��G�u\�f��|�*1|��vϘ��q��G��Epř,�-��j4(9���KiY���R�F̠F}(��%?WM��d�RV��c�2IBbt� �E)|������_z/-f,>[��:	�fr�_* �8���?Yc�2
��Vy��L�-��m��0U��\ElS��_x
��p�G�L��H��PI�#y���8�W�<z2P���e�y��!d����۴��,�].�ح����rf�#a��%�Ǔq;�x�;�^jM\Q�F����_��n^�����M�|
�4J�� u��`������*�U�heՠ�%B^Nb�w4x�f�*�]��c%�Z�uh���;Ֆ�Pgі&_��y�Z�({���~�m4^%7����Oߛ\v����%[Y!h���9���6'7H��v�dQ~�fWWu� �Yl�j�_G�t�֯��{z���`]���*�����Έ&yv6��sjl�J����w�uB����(�.;1<<f���H��÷�=�yU1)sy�T��/�
��g�씻�B����y��F��ü.���8j�h��Q�D+>�^?�T]��Nݟ#�Y�UU�V#��Z�,V�;��2<�:�"]"�����J{F��@�_�K��R��1��BH���(����IKZz��)��a�!�����>�$�Ld�g��-;E%�م��;�p8fs����7��C8��M�7.m��݊�h>,��"��=G�������������eM�8���I�p�P���Bm�ez���f̫.'��ө����+;�ʕ�qb,lT��N<��ݝN>��2������2����i��f�Ue���:s�zF����h�I$6�!ߓ +�5�Nq�\*C�=� ��������2��qq���(��ė�i�tLY��wN�li������k�앒�p^�0��WH)�xe
AM�P�R��5ܰ�o��t�a�M9��9�hI�\5�gw�(O2�ݱ���ſ+��?�6-�4;YO�a�7��W�@��6��&O'퀬 ��헺Vw�i$�6Kq9]#|�x6~��;N��b���l�jgtouY˯��S�"�X $2A��O��<�f��&�Ke�N���x)����I�:�H��M��3�_f�/�1j򻍒)�/.�U焋�ƭ�(l��n�R|�A�w$����}\�~����vOG<�6�cR��!�(��`�?���=���̨�u�c�^mz��i����Ei�Һv�Xr�`�tqW��x(�̾�f�SS0,H����kv���[j�CrG��֕�5Yk�9��E��Z1
�4�����f}��T�r:ԝz�=�B�}�F�]-�W."�e2��X�'}���׳�)�L�=��i�|��葍�,�Os;�̄�~�˺��z����A\��qI���[R�����&�c=������?6���jQծ��`�d���=�~>_e>8���W�!�� �;ХG��OBc�?S��|ԕEe��-3��I",�M�<����bU��8p��kB��6�R�	��A�&�ea@��"ۛ|�|��h��B@���1��_'�I-U�ý"��K�=497�Hu6�	��kh1��w��r�)`��x�����ͩ�Y�{�9b�D/��ƹ�/O6�Æ��h�9w��n|�6�H������v2*n��JХոD����d��W�\i��~�,�1`�
`�/���9�$ +���ٛ�-�r��cG��A��m��N$�b��:O����pv��������1F�|1)�\�s4�"�R'�?�c;}A۞o �z
�Q���G� �`��[Sh9��;y��\2�W\��^���=$E���s ��m6��J��6|k���
e�j�ǋ�Ef��Rh>O��T��>�x�I�`���l����e��lN����X�U��S=���_�=p��=ILu	{�fO�cc�߮��Qg�����xZ+� ��P�JD�)�,�ﯭ�4�d�Я^#����d��\���w�4I/�I%��6v�5��tl�+r�:���_c��}"A�qc,
Et�.[ZAa�M��5*DĲX}|�i̲�nm҈ZXr���F��� �ߞ�]Qr
����]"�!W���p���s<)��F6?H�dIV�̀�g�)5X&�	�~��?6qa�oh${ME��0��2���ߊ�z: �VZo�"���-V�/�1QOF%_��dy/Qix
�Rk?�������M��o7�4'=�P��������+ ��C%m�d
���=��2�a�J��G���h�N���v�M�5�n��+��z�U,g��~!
��J��r�R�P�-�9�@p�<�Wi��V�e��t�Z����:q��J�O��p�:ԨsZU�QL�YY�0��FZU��;7��+��XC�~�ƓgR�qybހ�l�U7�y��F��U�"����Z
�Eo�D��]��=���!�rЧ��@�%��f�V���#�PK-�d��>o~�uw�9�ۦו+bby#̔H�V�?��>�jR��s"2�Q�9d*9��ᕩ%�(���C�ѱ/rdB��M�G���V
��k!2&#���nv�R��0� i�3*x� ~jU&��栺��Vy4p�.�kV*A%ˢB͞�ң��VR��u`��>��׳�@��`A���񑲉��"A+��;������OmM�6j�0iZ�+��eBcW+�vB?���9f<��P	���mÒV/`ų#~�Z>5�(z��l�zV�$#�ŢY�Ҟо+≆��Acivħ�s�����P$/U�����|�M��L�>p�����FF��o���s��!n�B|�ڌ�)%�'2F����g6��j��/��@�lqg����ї��G���bC/� ޢC*i%�)>�ɋ*b�B|fx�0-O��Z�0��u�p��c��=��S���`0>����)	tzI�`�8����+a1M��<�(��()F-k5��ӌ�N��I��t���@�A���DQ��U��ě:���	��������`��L!��<�)�kV���v�2tb�'ADM�x�Q6� ��qH̆���&�4E^I��ޑ���YCP�l�����ט鑲�/��^#�c�-�lࠇ1��E��Sy�v��	�_rZYS��~3{BZ�E�põ�|�ͫ���6z�ښ}���R���*.ċ�ӯ���K<�oK-Ru���0����%���0��5{k�0���԰ �8%���.�;�j��q1/�<��(�p	N�jK#�9�N�Σ�BtU���/QP+d�xA�h?'oO���b��s�$�t&r�XUI[1A#4��_0s(��q��<%��3�aұT�Re�!��������&��D{�m��	����s@ �Q���d�@��B ���2������u�U[�|��D�|�ʨ3-2�Z��e�g8�
�/�eYl	��?%�%�<:U�+m_�pE���Me{���ߡ'�,�2 r��a���e���_�N^_�-�U7PK��I�q_^�N����˃b�'��#;Z�YrŒ�����2nk�x�� �p%�\׿�'@���/��r�@���B�I�=�ԭf}�i�ܸ��L����,-�l��}�����[�*�)i��+��8ܑ������Qz�R��vL����Y��]I�k�<��qRlɥ��Z�(�򳁯�;�^a1�l�� ��l�ބN�� 6�����/����x��w����9w���rڋ��9�gw�-��� �������M8����3�����8�Yjx�ı�����1	�
��� k ʨ�y5�/6ho�.�e��7o�ݒn��x���k;��fᥙ�_ƏO1h�I��X�xh[���|�P��y �)�Fp��b�d��˔���2X�yѹ@������ő��$�A�1��
�RC�ُ!�2��SB��u�&%���y'��5��9d����_�����E�=���z�]�D1K�q���`*��ZEM�ﲽ�-����}���ev����S�3��d{�۠>�Ѐ�/�?�j�V6�F�>{E\��笶�jK��{�`{[��x��w�(��!��w��Б�ܐ�˕�4�@H�6։���WJSZfK�m+V%%�}��<��#�7��5V��TRi�$�r ��1���>���06%D2W����o&^w�@��TZ^f��6�Ct�����������.���nC�,�6ۛ���J�1����;x~���2��Q�~xn{5%b]��l�6�H��+�Q-����U�iNW��-m)B����Hsx���������2� ��P�߲Ia4���Jͤ�MֶVE%s�MU�H:91ڦx9&1�U�?�H����dN��ƨ'>�R�4p��P5�F���rrD�����z���s�ɻ�QU��3� �B�qs\&����*�9��O���P�a�E&u�>v�_���@<�[���Ӳ�§8-*A&��d-�y�F�/�f�04aUP#� v*N>�lѣ}4���W���K�a~M ��;�&(̻�O���o_%|$�T8�":m_��[X}e�5��6�6�27���\�~��Mך?f�W�����o��Ȱj�f�۷����Ec��)>K��nJ;;�O���Kr�#t����zGB��^<�-1����vLSBD���_f�*�綕��|��gr%A��|��o'#�;�{Qyc�G�Yg�j�2ż��{��Yz��������:���P��>g<��Dؔ�R��Y�;�F�e4F�S-��J�~Z��ҴyBf��w&>Gy�}�^.�`�KͻC��$�"cI�y+��K�*��e�)̌
z�{DN�(q��#gw��H�F�dn�G/�wN;��i��~���T�*�5i,o�I�Չ�z�}�2�����@���wdҡT�y�{s�����3�$��Jl�2O庋[�=r����m%�n���>�k3���Ԍ�ļ��_B�"5�c�ׄwq8|���� m��TJ|��L��Ԋ�b�$~=�M�� pCV$yA�jS@UX���u[]��e�
*^�<(ܭ�/�aD�21Ǧ,�����<̺�׏\,�?=$��������!��͟_zJ5�T!�mfn�I�� �iD۔Ɣ�����,5De��>����x��񫶦�ᫎ���
$B�Hr,-"�$/釸\�4��g�?5�,�̷>i�z`���ڨ��%؞[��T���1���Q��hU�܍6�a;}ۛG�ܙ��4��]�D��Ĳo�.�:a�؀��H1���U�L�v �D�^	5�ѐV��OR�3G�=�_�wu5\�lvq��m������^3�w�D[��jT�;��R���~����O>.��H��;^
X�D�pQ!x�vk�&?C���;2Ҩ!2̓8
����H	{R�r�9:˒��rㆢ���irx�7F@����V�5�B��K��GT����H����3��!�ӓ�u�:�dt������M�-�C��@���ˊ�N;7m�-����t৽�fǫ�R*�n���2<�c^���f�eZ�,�ͼ5I�>2�и�=w0�'�@��M��)L{��H[�6�4��7��kk�Z�頻%$��'ϗ��{8�*AE4�o���m`�����>=,��D�Z!�B�J!�
a?r��L:*?���4�����V@\�|&7]LF�ԥ�i�t������/��F&��͠zԥ�C�u�"�Di#y/>��ja�7��ƶ�ͼ��!��՚�N��i俔�Ԛ�2�̵~/_e��M�;���,��S���n���XLm�`��Hl���۴�	��M�S���3�+���#�Pi%�vʀ7����T���{����R��:�ވ��6|��E���E�x���ZU8ľK;Ý����a����� <��a˲�"��h���Vd���I	�&n\�F�f���A ����~o&�NTEz�N���tD=�V���7U��~�֚��
@tv�Ԑ��-�`}��r3��wt�M3�?��fap�Go���9�T�Q�1i_V�i��j�`��xU7�E�e6Ҫ�w�����~���V� <~WYhq���V|4�Bэ�t,�@뿜��	��:~�$/e�|�y ��$cg25�*��fh��q���F�r���c�c�H^qh��:�%�_C�ݠ���^L�[�K]����%��O�?{����򥧳τ;GT����������&�< _���ګ�2�����r���zyF��.�U�j��2g�2�b)sc���jw�=v�n�fgyj?��E/��k�|o�ى5a�{�BS<�P~%b��6��J `S�o�Y�*�;�)�_e�` ��~8�a�(�ש�ri+fn�YB>Q"�ɖ��*;�Bx ~�I�<l��Eٺ5C��b�b���8?���q���i�{c��9A��R1G�Ɇ�4�P�;��LOey��j�5�l, T`��� ���}�S�?����¯�o6��5w!5��[��S{Cc<�W�&�L��q��΀^�`�3N�|�N�;�q����"�f%���pw�mw�b��-�W�i]'/�%^�鐉���oeۻ}���,8�<Z�~�*=pET��?����?!���b�˺,zip�T�ђ��ƀ�A<��RUQd��%��'�c������^���hAŬ�x$C�i*�Y.����U�ӎ���A��x�ܿ�^��1�X���6����O,���ͧ
~�������ۘPB	�19>2D�v+�?�]��"��$����[�B�=Kw)�̭�h�Iu��bhӭ��an�l�e]���؊�O]|����3�Jː�݆,O1�6<��;�k�=΁m|�j�㞗� ��}��t���a��Λ�T�-�E
�D\�oȉ���!R�d�E߉��%%?k�FF�tώa����f\Ow ����C��3E}<���Ww(�\B¾RJ��J*ؼ��G�XwE�"(flw>HF���1�Sx�V��t{JY�"���J*\exL��*Y�}���xf[�D�b�*��p&Ԇ�rV=[b���Y@	I���5)�[�h�$�����~�M˓$kՊv�m{(�	!�=���،�3q*(7V�l�Q��w;�N0����12-S�˫� R��ȫ�b�8/q���'�ċ��ҹKҽ��'�`�(�&��P��Q��N�*Ç4)\�(}2%V[�K��ԚtR����lq`�E�=J���<O����`�?,m�顠޳:�����y�mk�u�4%{����ae�꒛��Ǉ>�,��\�
�P#7��V�I�g��,�m7��0,>��C����߂W۬�/o�M��V�?�k�#��ó$��tyy�΃`kA22����ɡ�]8��q/��p)���o��D딼���dS���k�@����z�-�;�����W9s�� ߀6C^c��c;�z���_�̧��R����b�P9�	�#�`�L��n����Ĳ�����<��}�!8��6ٙ�)��[��cћ����qs���`#-փ�h��y�,��G�o�S,`���{$��Ǹ.��9�IV����!P�nR�y��e4v&UyR%��Z�6�U�}�m�K�DR�d�9��گ��Wq���b�����L���T[��E�yK�y�Ή��|5p��lU=�3eg�L֘��N�����՘UR�gR����e�6>7�1D��d[x]=�Rl).�|�@��<<06�mn�)���E�6�eg�V��X0��ȿB8�@�p���)�ĸ�{?���u�{��7Ԟ�nZ��F�d��uR�=� ���;������
��p��P�0M��Fk�6p�;k�j����������F������y7��I;�1����U��0g�:&]b�bu�� ��Hʟ�GR�sA5�9R#he�.˻��������:e�"�[ӣ%H�����E~���������韗���<!��z>�%�x��&�
�؅-�A��%���Md�j�1��m\S�R�eR�=�ͤ:-�q�Ȣ�9�E �J���9_�/{��`���,Q�\���c��l��V�]��je��r��D.�l .��9�)�-���5A�{�c�����&��qa	���vk�D��,h��dmx�zፈƸ}��	?���8��I�ά����%Y�$�j�B���7ωoڀPz�;���,B��a�{�U"B�C�A\�C�Y=g�tBj]l\�^��ܬ�[T(��S�NBձ� ���$�"Wz�'��/�[I����/�VJ-Y��.��!x�Nw���؏�U�N��?��`���noX� yT� ���/�����-$�� Ļ ��m| �����H�kQ"���9�|���u#����Ib�]�^Sv���s��4���FdT�u,(b�
��F�YC�':���xiS��-���~�8�lEZ�Dĕ��?�u���?෈���e_��8��k��s+����n� �<��c�yoJ��"[�[ݯ��Y���u苫�2QJ�>i���k�_�'p�5KK�����)���{e9'�] �.�6'vl0[��X�Q�BLkDW)�l�g�<�����K<s8S�R��Bp��%G{��I�E����,�:�1_"/��oY���(�(cXV���~��]-͸�A6��8�.h�8�;��%߬LM�]�T��ײ2�U�{Y<�aEB;,\�����ro��|K���R�[��k�cKq�������t)����A�WjU����ݹ�!V`8���/�RQh�]�I�I.�����������"6�x�c!����XMAm����f0R���S��_Zؽ8���<��1�閁��Q�5�K�ף�v6����WkE�xL�ZӬ��1̍��K,�L�ˇ�_Q�)p�m�n��k�֋�P�jI!B�fs*��R:f����>��潉�(�p���[q�ui���;��%��)�ۇʹ�v�V$��c��RXc23���֓L�W�%���2R����%�����|C�
��4�;q3���D'+T�^Ź_g"<;F�4;�C�1��\ֿ{�3S���QV����_1���]����I�D6�Ԭ�׽nȓhɲ��0�28��׃�)m?�"�6�<��BSN��g���n��/�#=����a7�`Ӛ�~��~L�{�X6�A�:�\�ԎlV�= &�-��"�KO*����Ap��{����=��1�����8����4�}X0� }����(�m�Q(�ȁ����c]ϑ{0��
{��H���a��gi������`R�q�DpJR�Q��צ�_������T~��k9#�P�X���B����I���U����Gcc��R�T+�	��;�]j�,�K��v�m�A5P�5/���Z�t�9�Ob㎔6L��Ga6��ܼ��L�7'd��ԙ��©`��4C*�	4��э�U������;�Q/?��(K�Y;�M���8���ɋ�����j],!Dm���'S�el2	� �<_�[=ȅ�Z��ԍ��Vb�8�e�2*����^X�ή��ƶ�R�CCN�3z��2��η^�ܠ�ׁ�T�i��H�{^(�v��Dxl����`�U��)fT���&�qOpRc%�M�H-a��o�P�X1���?�np�	wǓ�#���4�#��˓�d7UܵE]�΋�'��"V
U/��Ѫ~�o��Q���Y�M���~�+�A<�����'I��z-�%V�n���"'�����W@y��N'T�̡8�l��>	'-�P�{D���_:�7u�N5&#�询f�2Vq1��~��㖖�Hj;_9�i��ٿ�)������9i�o��H�5D�����������5>8`&�Xr;h5���$h���+2���`���[@��\�ȏ�[-��N�מ�'�|vG�u�iWZl��?�¨��Q$�l�\�� n�W1��	:	_��I���X����}�b��l�C9��m&{;X=㈮�@���!�#��3kmB8>.F�YI��|��,�(❙5+f`!eߧ�%�����B�Yh���B�U�<P�u���`�ˀ��=\uM�GN^ʚx9�e<�4�߀:h�ג.P�]#-`�;��?[��4"��'�6��v�ތOӰL$H��csz���-j��Ȧ��y�<�~����L��)�}��1����:rU�S�B۲��a�g���N��z���C�&-��<��{xmG�#�\?��43�".Dl�B���S���o̭`���vC=��`��X�p{����� W�"��u��i@���4u���pD�M��;Xv�ɀLv&�u�J��n-�����I�)墷�D��=���X�W�;gٞ[iCB�k��^��䝧��������8{�.'<� �U��W>�R��d8����E�Oە�\���qd҆�a�yTT޺�4lI���BI��"�!�~ˌ��'5řfx�0$���YH���Y�p��!Ls��?o�%�|8L�{Bx�T�����+7e�k6c�j� T�r��)x7o�FJв}��(�2���w4�q�	�<-��g;�+�@(�S�ʿH%ʵHbCU#)kv=��
7x�k�p+*p�1����L�( �b�Gy�aMAOM��Q�$~&,ݪ%��=���l�@�b #^��]��9�7�gʸ�ڝY���-z}Pk�Co]/����hj�bjU`^�p�dA�.~������S�a=�f	@����ׂM_P�>
3���t�)xP�i��+V�(�8��f(�{��^�
I����$!Oϣ �[:�LT��lKZǈ��
��F؁�윓LM"e�w��/+��}Qy��WqPm�p�������|���E�>� #�b�R�	G��Y�3�e�����|��Z<o�-:�O��B��In��[2@��	��8���4f�_s�J�����ϲL��]=h:�v*���,��[�{�b3e�Aσ�%pf��$Ȳg�A+���ϝ�x���6I2� ���:��oJs1r�1�d�7N$ȇ]7Kd�I���#�����:7�ss�Z3�\A��{2	n�Ǌ]�XA�{����}���o�S��2
�q�{���S��5p�  �o�JH"� טE�B�c�5-�ϣ��L��=�4��1����{�c�-9j�u�� �G+G��n%-K����ޒl�i�,���C�J(�@g����^'8�'퀎�Z�$B�Czf= ���V��&e���|D
�}�0"R(����H�~���I7=��R�/Mş����U5qS����p>,�4ĉ`���״�O+m.r�z���j�n΅��-��iQy (��Q
X*��p�f�����ğDV˦�#6�j�e,5�{��AP*?�8�\��0f�j����!MO�|@ ��;�$�E�����{�a'֮�
�EIa?��C�R!uw��I�w,t=O�"��zcԹ��뢛�gH�\-9�,2��#Y�VD����������?��~�gj]5�X�ԼQ���j�L�&�-�h���*��e�gb�A��+���k�nC.o��Pݑf1)ew��g��N�ȆȚ�������L���1n29��\�A��_M�ȃ3j�S�i�:�� o�'y�J���� LO��8F��{�	xX<�1%`��[ E�±-{3w��-<�Q%E]��$��
g���$~��yH�g�_�J�e��[׽a���@�F�8�V��K��-�G�q��'*?���#r�3q1�^=����N������|��XQ�y ������*MG������F14C}��w�H{�a.n6y�*]&��P�ZZNJ�����VHY�
��)�`����������� ���fד�YL�!��of@m�#���K�[-�z��@�������~f	�4���h��=f�V[�ِU�����#m�R/��f ���w�Y�>�VOuHO���&&<3�z�Hr䏹@9��t pmڥ����t[#p��nV�L�Ϊ���ɛ��gH��:���V�c��ki%�}��V)L�Aȩ���r����*qV���<Yg3Z�	]�,nl�G`���(�OA���@�]�vL��Ђ����'�Z@ ��ۇ��+�t�Uʩ��/'��@��~1�]�N΂�~0. �+^<[Z���?��躊���2W�T���F�^�wR����ۉA�Mֆ.��"c�-���i0'�P�Y�-�a�]W�tXu��8]U���P���ص�s��u���k�r)�d��[�5�7��U��J�^d�ok�lP�]
�_xl� U4g=O�7I��L�2�U�Ga��XR��?~�S���B�#~��YA��ht.h��P�F�\���� ��VQ>�.�Ȭ���z^�rEy��6gV�Ϭ�V�w�ĉ�bؽ%�Xi�*C�f9r0��9Un�l5�i�E�������s�N ;Q���_�zW�f#M��S������	�*?��0c�|�n�C�K	R�(��|����^T�XڹP-�|n�?d���u� �+}��_�0\�T�U�h-�!��������_s~[3�������er))γ*࢛g��f�D�"\-,�/�tP>�Y��<H�
�q�`��]�k�1�� �O�J��n^�'���2b���\`I5O�Z�B�N��&��n5�Z����p�ɉ���(��-��b	�Nݕ����+�W��<澈;�,W��P�"4 ��F�\a�y�N֥w��ϲ*>��Ɋ� ����S�6|RS�,�w�V�_���Eֲ"C5pdH�_m.P�J�W0����>%X�6�Q��b�Jt�0�%.�b����	�se���6QlK=OU�z*5m�/(JuSsĔ̩ݰ{���j�6$�`l�a$Z�Y��4񋨠�G��r�lW�B�@�r��E�w��b��1�TV+��3Ń��3_ǫ��%�?��`wE�-e�Ar����*`�
�^�N�H��G�t�ƭ�)�|��L��\�4X��(j�=%�`=�8*�v4+���6F�ZF�|pHu��ڀ��d����|����_wH�a>��8&�ե.�Q%��9���07?B��;�|�7W#�@V���Is�� s��L	��.d�Q����Q����HC� ��M?���E��_�ߚ|����	c�!LU�ǡ��P�V�_�y���Fc�v줪eU�c0Y�G;'N�#t�]t�����M�7Z�N������R�������A�8G۟��I�Z�]ۀvTB�
̝�=bp�Z��7�_��VGuZ[8����c�C��C��v���<}:�KQ��2Vv�R�'w���47J%dSVc"'�3,0r�.FZȀ�S,Ј8�!�N�NY�Ya��t�,<���-i
S��}�0<����/!r���J�ck���/1���q'20ҡ�\x�|0	�*�'����,f8�A,raN��"�@��W=�/s1�G�`#�9!<9�nsS�5Ħ�I�ˑ*QX	�����u���Ч1(� �pk��۶����Q!c��\��}�/�'j�/�d��|���-�$��P����,�U�)Ӷ��kd
���B�B���8�{�_�����P�v�t�֝k!��Bʅ.��v�Ũ8GQ )��
��%�p�%�*��F�̖=���O� �����^�Cl����w*1uJ���I�UA5��xا'��t��t�bs�!W�M5�\�R>W��=��V [����%���H
y��N"�ҧ���ۥ����+	��8�i\T�e* ��H���1 �\X�*�k��J��(:���iΆ���e�bI0�-��:H�����.���,M�
�b�}�/
=� �e�������~D��8�21���Q���f�u>M���*�n��V�8�����2�ܝ\������m���,M2e��U�CA��P��l���ø�="� �#]y�ŉ�Ñr�/�ǁq�n]�Ԫ�q%鲎l�#g!��-(�� m$) �SD�z�q��bUr�u'���Rt7�7���p��
	hJ'��`Wb��sb���ZmV�u����Ϛ��6.�t#B���w��N�gc���7B��)��]R�a��UZ���p���l�>�q��Tdq\�?N��u%����>���z��Y�D7��F~��J/!�jW~�(��:�e���X%Qǖ[WL� f�`�lyf~��D�(H$�Ʊ��*�!�%"��i- ��w�=hW�ׂ��:<����r�5�����O۪�pX���3�|��b�^ �Q%m'!�K)mG>�s���
��C���Ǖm�J�⤼�懰>�O�����HX	p����.hH�a��6�H�gH���K�Z�EC�P�o���Z����j;@�',Mt��?�^����ū^����L��O�b�'ӶD}v(h�;s4��D�h�,5�h�l�!��ju��}CQ�.�Im��qY��)�����Y�I��Jn������n���u��G�v9s�����R�Uw�%�����FV�v����7K65�+f�V}��&�I�K����E�^KS��Rh�z1�����i<�N'��>�?�6 |ƚ��H����=n����G��f�?�;�ߨ��æ�LzA	�f�d�}�Z٘�Z�LSS�	j��S����0Ç�����L5�0l2l���hFB�>�Sq�z
9w��N�}�z�M�N�
��|ډ��?���%�,�~)8��>�T�(�w]5",�_$�|�QW!�P3�VG[��+���Q<�!FR-��r�I��(�@��\I7���hg�=<k�^�c��i#o�b��sZ��W��H�Lu�Ù㌫�������}f������~����S懆|0�F[&?����6�]3�R�0`��}8��@��_y>��������R0:��m�~����/,�k,a\�.P7�|����C~s��1���:�"������ty'���	�@�}ʆ���|�S�xQF��s�쀴�����+=PL肋�����d�i����j&H����\�����H$n�e�L�n.�ׄ�`)��. ����st����T5�Y(��v�<�IA7T]$~b�R��{K�_.^��p^z-	���x�*�'�C=���|��bN`��E�U/�bM��؍r��RV9�e��3ف����pa3����=���Sc������Fq��	DFP�*CO�o)�.���w����$�����7��[б{8縋yZA��&B7�}�Y�Oo����5F哞���F7��-8�Bt���A�#�N���O��^�䀐;q�>ʩ�ȅ�I&�Jڣv�vq�����-��rS��>1�S���bQN�Vh����Ѭ����졠�d]gE���q�~l؈=�iK�a�i�˝q����]u*k��\Q����+��O��O�[��l�pw|��X�����
�m��P;�4����c�*I�Oi앑T�2��£�����v�4���7�GB�<���R�"Ʃ�z9��_�����W	�$y�ë�j���^����Q:^�W�5��3*|ǴE��hĝ��)�`:��۩�+3��QiI��4J[��zdߖ
�\$�M)��IT�^�]r~V��(�ݱ�J$6ߍ]��&)����iy�?!5g���U}@�tanR���Vaۤ>l����h�0#H)xѱ�Ant��G��(��8��@�?�CW���0^L��\�ge�pymN��-f�-��K�"VT�c$�s�p�X�w==	�����Q����؉�U�W%2KL����|�����9Y���f���L��M��p�_�j�4�k�w~����5��`q��9�r^U!'�������Y3L/f�&�52���hr�ҥ��*p�L6�,��z�2%
�H���W�VZ��pm	�Ɖ�j�{�W@S�2�)á>���%)V>��V��k���e7 TG���n�X��j�ժ���;Ε����d$��@] ���n����t��βP�eSϟU�0��IA`�YQ1bŗ���5{G��g)�5�!A��cod� ͦ����Q�qf�Oߣ������4-ġ<��
E^Xc���O�8�BO
��)���b�Ҽ-��x��x��c�Ģ���SnCՊH��Ӟs��Oz
�l�8�����a^���`n�b����~�X�9��M���'���>�l�����w+�	�oZǫJ T~ƳN�� q��@����A?���W��M	�g��^��,��6�\�'TF�XĂ���q����碊zR�U~��e�3�p�&�5'��) WI����R�a�xZ�m���b�<��(>|3\���0sC�	
��Q�D��+�X���aV�~���pUQ�kj)�bE�R��sP\8�L���+Wc�S�
���# �5En�Kq%�9e�9��#͖���:\Z�eOxJ:0ɩW�N���GM2;;�cdk���Q����4�� ��
�t',�1=Wz������4٣�@&m>��	�s����pڊ�~ o�wʤ`@�����i��|T�p����/\���Ƅ�y5An&x���F�(��?��=dE����L!6��l�3:\�d��jD���n���ͩ$<�(HwQ|������}�
怒48�o�eh#���s�_qn���P��4nUV{�T!r1~���S�K��䛍iҽ:�\����Q�L
��@�;ح_����~�X O+��п(�|3휥@�I��+Rq�.�=2$n�����;������0r7ٚ�UL�b��Fl4[2��U�>�z����~N�X�z�@�"%NAZFiH#yPH�^���G�D@����h�9��dw�6�ٿ��:)+UQ�A��%>�4F����m:(S)�����C �]�)��sv,���n�2/��L�����:��^�C��3��*R+�'��mz�↛_b8�1W�]IT�勵��8���]$�����&���ڱl�m���Q%���@�s�C��{%r�Mf�u�i�x����M�d�����Ú��%�a�7�����l껞%7�A{����U����-�+P6 ���Z�1��46�9�����EG��-��ܲY90�\Ŀ�̩]��^�mJbh�̐�fO���@_z���ih%�N!T��~d%o��P6�}�!+/r���TU]Y �9�Mb���
dB"���9y%�A��|�� a��٥���QO�����U�[�w-c�w��G�,6^.;aŋ�ϓ�?Xt�N�9K�X��������)�o/P�*��$�l8Q���(����4.w�;�c-�������������7�}����t=�
�����{Dk��G��_�G�"rnJ���nB�����0��,�/XȤ],�<�D���
I�g�N����K�3ҳ���Q2�M���6][��0_��3�a���C�S�iP��&)?�J���n ������b:�#c�Q#��2��,���2�E��j�b���V�|���'ê�����9 �����d�z,��Ʒl�����#�����Ayri�%EU��\|Waf/W(�����vω���)��)ϖ�t�=�K�y�M�^-����ܲB�	XM6 B>��U�.��79���a��'�Pr��q>-DO��3�5�o#��ĸK�������b�����K������J���J[yc18D�	����S�o?�]=��1� ˿��l��ݦ�uߤ��.�����˅�����ڻ��|�L@��5(y��R�����n��yFi�u�-�쁒�K�m�� �lW��d�����%��_�Q�+y�1]�1Xf'�sf�:S���^�^�$#��9��@'�,gޜs����١=�ח���CCP�[SO�:u]���S�9P���Z��fg~ˈ��O��/���z�MW�adw��'�r1��w<�m��&�'�#\�tWYW{���i���.A�Z:B ������Nw��⟨�K�2��~�:6V��N����M6�b^�+Ǉ��üN^Զ ���u��r5� rp�I����s�χT��t�t��e=Vj�G{=�N��ˀۇ��ɚ������%������O��.��Q�_�{CK��w4�������챽�2��@�%��?X׽}�i>e
`U�]z:��5�I� +>t揈�xO��^���>6��O�������1�Kϧ^�|�bLYx�3����o�i�h"M�{	���(��v���y~rRF^�"����MR�K��&%���-rI�0�ڊ�S�p;���}�����5�E����"o�8���%��bXC�D���(HOl�G��oI�$H�1d��`�=B;��3i�������buƯ 4h�������Q�
�p�`Mu�8֞��q��'"\/[�,�@�[��X�d�$��u-i�'E�޳[� (F���D}��H�2���Y#�F�y�o�'4�H���p)���PH�,tʦH�H����Y��M�3ړ*��+���{��<�ȩ�{�CV�j������Hqô_*Cڒ���/ zy��ݶ�^�����L�P�j���n�3�5���S��p�)��+/:��Rp�-��;j�������>Qi=�'��;�y򑛿s��M>����7�I���#�p�/�y8����7�8-�bZ�H�,%?���j����͞&���i\ T/�̍�Y��,|M��h*!�������_���u&?L7q��2ī�eA�^~�j^���'��-I�mL�{}�q
D��Nk�ZU��rQmM�
�g� �.�k�5�ﾦL�k˕�y�@��;�	5V�}��4�W��O��<=��䳧v����ɂ�ޱ�.����e��������?�B�z&�I��x�3���D2���GOʡ��wS�N�?�%�H�������<�ҌY��$�[#�'��E���#i����L	�`#�������_UH�DJ�CXN	���¬P-ŮJ�?�����W(n�^K��ƽ�f�^�����e�G׉�E���)�gL<���0Bi�6%<,̏:��qI��eU���~��r5���Ѻ��"S�ռ��ā�݀���S��C�����'��t2���@��uə��"��5/�EP����'�S��?y���qқ�W���#_��Qԫ�quJ矏���[EE��,4�}���^�uz .�(8*�8lK
�M�:,_�U\[?2 ��[��Nk�k�4��Jw�bH(}5B�f���Q�Wuѯ|ߢ::�b��ɡ�[�&d�i,B?}�E}���4g�Ϫ���������������Y�W6��o�l�����BgFȇk)Г������B+&���k�%M���h<]Q��_|����o
�cJ>I<�~�v��
�j�u�"^ p����Ck<M�Wq-ʃ�T{W�-��d�'�tl,|+��:ª�7u[�ԚP�+�z3\��j�6�r1ղР��x�H�T@�՟2���@̢X���}�+�����[�Tƌ�1���g�����BŻ�tW"O6�X��fuP��P�Z,S��z�/��j��k}�Ȫr��W�WѸ����C�'ܨ=璫.ZjΦ�-<Q:ɾ���]��]��_7�T���nt�<;��0�.��j��6[��0l�N�Q}o��[9�Zb�s	S9V�p���F�w�g'`0wWb&v��V�?�}��u_�j:��F��]�r�<�P�����ŝ�L�1^��7�7��XE�R8E���WI-��Coǚo�p�=g� �O>�XW�����ڬz��O������Z��Q9I��+���1���ŉvjʒZ�
�ߴ���c�\;5�����u�=6z�y��ٛF��=~[:7��^�K��x�p�m'�y���u�d/p{,��br�	s��!�;�R��1��c��v|��?�mO�	�2��Gd��ϼY�ף���h��%47�L�o��m�a	���ʇ��D�|�a,vx���m��W[���d���j�?w�P"}sXqI�e9��쯍�WBɁ�eH ����� �U����]7��}�X��^w�;F�'�Y���i쨿,��v�������^oٹz��>����&Y�m��t��Ie�����wK��H�_w�Q���87)�wz$�r\_���8�D�%S}lj��_n�u~���q�܍4unH%�Yע�Z�4Դ�@��F�nǅ`�ӟ�1��,�,��,�v��B�z�A�LS0�yqt���o'&�Yժ�9Y�o.j�:��妞"N��lH�o�����/A��n��b���%Ii��Ԥ��i�x�fL�6a���E�Dj���jTH����"��7�u�MP�Mj蔊92ێ,�&�I�]�:?Yطw폼�v��n:���=����<��@�<
J�8	C�&�bB!z�t�JE�ߺ5���}����L��(�H����I	��I��������K�6ו:	f̈́�<�K�j#5B1��4������"��$��)9�_�s)�����IL eY
3�=:�dym��r㓬�O������J�}g�r�ȈA��@�@�KRQ��谑L���O.Yq�S���mש�O��"�
_��#�?�Ŵ��r%[���Ʈ�}�gz0�N'�jŊ�WW_<��_�9�,�0
��vF��=��P�c+��ܡW��8��S����*:	V��u5��~��{�o�?�m�˵m߄Hk6{�@Ї!���WK*�Q!ɖ� �pC_R}� ���#����%�&C���Sڶ�9�#��)�����-.ر���ҁ��ߜ���"h�����	�y��������p�$�$�(%�?�f��g@�]y����v�>R���O�|d�5�-�u��/��E	��È�:���a��l�6�F�b 2�T�H6Ac�9����|���=��s�a����z�y�pdc)i�5��� ��Kk��Q�������I�q;���3�LX��w�K�$~JݜÊt��"��V�pg�i�GR�����0��տ��i���-h�I��HXչRd���KJ�!��@r��7'Q��E��BKb�3���ؓ��U'4C�~o������=J"��2��/i��=�F0��B �N�ݭoi���"c���3D^û|���d�L�b4������X��Lk��+mYv�/����Z��JD���c-����Y��-�@�N�v��ɦ&ɳc|ۆ���{'r�*�n����[�*M,���!C~ ��nZ��Z�^�~�\o��1�V)�h�N��˹0���a�	.3̏�M|�;��:1��*:��D�����&\�Ѵ���#h1F5S[��CQDn3 �z��:{�� ��i��)��L�����]�Q���..˪�R�S"P57*PuL����or���Kj��>��L�*Y_����ӥ
a��f��uNtU�Is'��.��9�em�c=`�����u���z$��W�&f��� ����n�D�t��m�,^���o���ЋM��I#�H��4���:me�bKgM�o�c��N�r��j9�����0�g���Z�-�����͹��q�@���O�L��) W<?N>��^%
��?�����g*�=Tꀇ3�!�#lV�9��:�Kd��V��.�¼�t�C�\v"��=�@�m3l�S���S���1�;���]h&�oa���ao.�=0���t��O�$�ߪ��b6{��˂9���u����qCd ����ږ��O�LY�R&��{� :�
a�D��:&m�������71Z�Wq�D3�r���@q��S^��.��[U�%�s�ڛ��v;xeJ��g�%��X���Y�l��g�0d�������#iۀ9Ϭ�����=8���E��S*G�M;IV��'��������������!n�9w�Y@?uο�L��8���[�q�ޓ���;����.��ſ]���rt���<��z��KS����}���=p��S������3Vz���P�'AP�0�0!�PV�/ơ���?ݖ��T���0/�͵<�ZdBLw���uU����`xc,��p�Ï�既���}2��a�[X�g��c��c)��d(;�[��`j�a�x��@)�mH�Ҕ�=��M��M1��;��U�I���cUd�5�
��J�N(Z���1VrP�+e?���}w�e{+�������FΤ
b�����ɷ�	�z�h�����E����:����3ܮh����Xi�qx���_U�MF�������F5;�D�M\X�⼝ml`�Y�mV�>X 4̩��C�IL�PZL�.!����rq�Z.��;2��vK�\��b�3���o�m
�}Y�B}��Br��9m�A��ً�J]L~|0��AѳG԰��ں���(����!�Z۰+OIv�����0XW~���ݥFi>W߰��d�i]�RHp��ל�TB^�� ��΀T5wo6�����J�KT#�F���.n
b���ρlr/�A��o�3?l�"T��9�&.����k���m�98����(���H*�?����G����r�X�q�N�h�y{#��@��ox߈�����K�`�V�}��05"����p���hWL �rx�OԌ�ib�Ò'��-@�<?���w#��)����oҴ2�����/ӟ/��XhF�sv�<� �}} c��B�S�]F��K�g[������^!�/�����x�k�<��o���j+�A�|j�B��'.DQ� I8�Y[�@+�;���#�����3�q_f>��
���uQ-��}���fW��Q=�����j��G�.�������a k���宼��l����]*����T�ۃp����[�$�0`A�%)rZz�m�/t_)�\�g�V���	�+���!�-���΋݆�Ƴnx�j��c~�&�̸�-єG�g�1�|��jy�Ɂ��"�gx�4�O�^�}�nOz�н�c
"Gnt��q��S3���7���H��`�	>!�p��FWX���O���j9�P�[�F�a�&`u���٬��zҫ΃� �Q�}u�~+}��H��۟�>���ؓD������56(3e��-?�}�a(��S%�ܭf��V��$% �-<�x֛j��?l��uυ�Ƕ՟b��Q�LU��"�A�>�-�H�V~��f���벉�'�a;6�Bj��X�mu�n��������A lo8��D$���D�Z}W�
8'b����+�* ��b�Gk\��}���L]`�x�9?_�b��YJ"hz�A���!?	(��v��]=3ņ�QA��]V�./�#�+���7�!@w��1Yq�m��ï����}�MmK�rZC5lפP _�
��ŝA��)��υ���'�[�2�8�c�֕��6��xd�\#�	0�-u�M�r ��}���;��(D�����G��sc����!�S�b\�)M���!�=)m��S��	�Mm��~pOu�����2���ȫ\eH��۔���:qƺ�"|�kl	A~ϛ�.�g�� ���8��r�@h�"�1��]���p8���z2"��GLs/n��%����Tx`�}�-�u_��؇�X�90���%	-�Ocq���R�pj�'����&F�a}�5��.�̯��H�k�4O߱�]�<v~���UNlA�<y�#�|��VLL9���i��fٱʊ���?le�ދ$�,��{��y�Z�a�^o�]�lM�Y��_�k2_��L�N#�����٤�Y?���&����"F�l��@�?s�����>����}�O޳+vߴ�_���(\*C�( D���:�����=)8a��k�U�;��u��nI�[�JӽQF�UX��Y������ٳq @�q:B�꿤?�9s4``5W��ɋ��^��n��7���,�
�/@��),a���_(�x8�3��7��3�	���  GJc/�I���� D¹� �"�D�8�E!��%����u��mrҠ0I{>+X�fv(a&#p]k�a�\�E/����o�Z�i����;T  ]�h�!�"��K���l� �5V\fmp�u�Dqg]�crs����A3�\���-](g�;&�Q�7{b�����I�
����7�Vc���,{�֪d�7��S+$��/���3Ҽ~�nM;���]n���bh�±��Pew$ˁ�]��S�Z� n4�^�G�6?�v�C��b�eFd�Q����dO�k4�M
N&]A�;�(���F_ۑ�p�J
%����v:H��ˤv�m���IJptb���5���<ܘWo��r�]�N�>;�.��k�<<�W����i��z������G��z�)_�E��^��Ӆ�:�!4����r�ѽ?�<g�﷞����4bHY 1��k�Ab��!���@-���L�^�0`',���x���ת �Y�t�&�v�"z�s��oT�?ۖcu����Bv)�Dʎ�����l7���j�"��"�>v�{��v��$�h?�4<y��@���=��]_�����8��/.�(�1V-p1��/e�_��y�����,����.��M2*Q)��l�鄆�G�ݷ�� x/���5�3K�[-za��rQ��Q'-R湯=h����R��s�6�Y��"	�/�����y�Y�@���*�h1���	_���r�Y�}����t}B�+rc����\�� �)fG�Y����{l@����U�w�KYC�i��c�z����H���gu�ש�z-�&`A⤈����~2�]��ޫ�
o����U�x?Q��֦���t~>�sS �ݺ�֩Mfޕ�nB��3�"�\&��-�C��)����rXβ�?���4�`��hE_8�iܷ:{iţ���BO#�M�2Y@8'�J��Ȇ4iVw,:CC�4����2�emq_fM�C�K?.܁��s������;���$lOC J:��6�bf���/d||��\
�Q�~v�g�]�ڰ~J�E�+��?����~ߗ�2߿������^���3@:���i�M@���&e����()��/ӗ] &������`g��%u�v����׋�#�}
��>�cз�h��"I#�� "���[��$���Q�(t���	>&��B�F{�!9����)r����Fwͳi���{7�/�]�YU4.��=o^b����XfYD��"�!�U��I�y)U���܎D�mvEV�-�%��������f�f�ʕ�/�����6��^VN�N�m�,T>ށ��+l�geЦ��;z0J5��%��Ŝ"��u�� lȄL��ϲ�A	2�yK&`�e���5Y]�����f{���/S�m8�Q�&�Wo���3�#��Ծ֎�6��������/�au�g!��P�3&0�B|�i��dGF茖��6Y��R���R����XY�=d���~X�['�+2ϳ�/mw���X���=}�����a�8�I��V�p��g�P��}b��p�xf$���od{���h�ѺF�&�{������0o3�B�sgh�<�*�3AhNK?�0��4҉k&%­�7?D��>�τ��K*�e|gO%.M��y�"��+��������x%�^����7��4^m��k\��	��Qœ�lH��� �5e�܆=��I��⒔��y��7�l�Hr*�!�@k��܎��j��|��x��x S)}nn7:���`��e�q(Vl�u4�V��n���&�a��π�ީ
?��]�)�K{�/���U@�g j˪)}��T��@9��[���ET8;)�Gr+{�(�t�"}�'d�13}�{O:�ñ!;~�~�~�y;��{x��<^���s�H����%]}t�Ѡ1)�&X�%��0J�=;�f���V��L�<�䯗}x-lx7s��/�oқ�&.βԾ����P@Շ��b3��\�UL��g�r� ���V(���,Ƀ=����P�fM{�5�E6E!Z���Tv#�g ]�V��S��ˬ�dH��MBn�|d�	���B�8��u�rJ0��y����$�q�[�z�8�K�K��oF���<em�Y����׾~8Iy�kQ�3���٘aV��i�k�D��X|y�b�����A�/��J�Ys���[�+\-���K'G4;����#�af�s�aD;��|A0(j�̏bf&-�<��d��
�+aTԜ*�GLB��8
��cb�R�.yI�ăo�h)^��,}�֭'�B\��d躷��ס�}x�al��7D�kF�_�S
�\����N�Rs��JP<�B/�`><a�4�d3��w��� }.HL���NeOu��,�Y?�!?�*1��48oxzA�����V�g:�\���/����@�7u�6kh����Z$>2���]ԟ:f���ڽӳ3���pU�a�F����~��z��:�� ���|G	�ߓN_��������Z���J��/�n�	߀�p/���:r�y�BJ���v^k4�	��H �2{��!P�����-X���(
2���3V�Ʊ,}���h�=�X����C-h� Æ�Y=����B���/`��$ϫ�����f7~OE��nn"f�M�7fI9jb�F,�@������ ���z'�k��Ef���x
��a�=N[��;��7�Sw+�Lg�JNߌ��Sh��x#����;���A��}�{h��P��3b$E�v��jK1>�6����c� �zi5@���N�
��}���)���ݓr������-kͿ�ป�o�䧀B6ۢ�	P����}1�rX�?��%�]Ī^�d��׮Kk BTw]���g鐦��+��C�UB�_о2����p1^@22&z׆����S+�udK���и����[͗�=0�5�Jk�&}� �v�u�/���}|N"��p�Z�A�P��s���M��% ����4[������@No�f�@��=}96�%a&r,l4��� 8 <���r��۵��|�";�qP��)�a�����`j��f؀CtO� ,�- ٌ��6S���H���:`ڏ�T��^��gT��M������/��&'�D���}x��҄U�����1N,4��lUZ��%C������*E��P��]ԃ�4�ۇ\�t�K���~1w�`�t�~�Gt%��r�`�8Y���.ٖ������3'�<Q��S7��7� K�Vo��D�N���a~�6D��?8t��N�{٣߃�����>�?��ya�J~N�Ψ���0e����j���?��)��@Z���f��-O ���#*�MH���z������@m��r��;lёpq'�<B�7#��>�iy����XȻ����r��qm%�K�j@m����y���'=��u���ŷ�^h���y�%<��ѿ(%P�t�K1]g��ʾj[HZ���`w�X�j�)x�%A.����e�TOJ�ˁEL�[\���Te�v�ޯ}'�]�������[��<C�Yw����H	@�K�X��^p5���w_���e~��K�.�����K�Y�ܻO��m�g[L����,CqZ��A�N���0'�9Ogz`eF��.�}ڼ��{ݹ���G8D<"����C��>P���j�^�jPjR���ޛ��\(]�T�w�]�������u��|JAXm� -�u�6��?B}6�䐊ˠK��A����\a%:�Z��o�������H�L�DVW��][ňw ����I$k���y���hsc|����f,�;�+l
��"	�.����}�B�eXǱ�����_ ��mպ\Q�K�o�6Uy���P�P�ͤwCA���]���.�ey�e��K��`�=^1�+��,u��M�zF@K��̇��?�7KS-���'�݂�I�B(��h�ڐ�*���x!*1{�OIG
Nk>�8Q"Δ	���ÈR�h5˗8V-{�rT����V[�"BZ�:��"�@O�K;�3vC<�8@y;i�q�����6�$ �߉��U������tW�C�H��5�	��$����-{��K�t��1���.�+g��(��$w�=)��Խ���P�~���Ls}��' ��10�*��L��!;w�FD��}��:��5����1y���d��ƱmJ�3M�U5���$B�tv�5[��܀��&��٧����F��&�!��0{S�nX��7�"}�\� Y!��?�j%�ˇ<�z:C�j�=��oQ)������e�]��{^ ��	�IQ���	��������(��u�����8���ii�hh-rT� oq�*	�Ɲ�����<�iv,�}3W���{�lQ.IQSʭ��+_����|	d�u�YbQ��?���x�s�NV���7v�x�X9a�=���g����le�ۉ�}��5��@'C�o�U7g@�ct7�w�Ksp�B�sN]'�$`q'��0|p�I��n6u�Z����]`��Zy�U�v#�9z�uߪ �[�E��fQ�6��|Ic��Z'�� B�\(ӭV�m�깩���'ڍ$�Nĕb_���X�.p�x���O坮���������;�	O�Es]�L�{�.��ٮ�8t�w����Rz�FV��K��t���1.r������u�H�1n���2����v�f�Ć87�����V(��َ*vsρ��k5�d�j���Z���%a֯no;��3g�>y��*�4Wt���=�1%4!;�m�e��ws�![�3y��'[��.��p*�O:s;��WT8�����i�ŀK���GV���Xz����R����<�'���8�^pp��a��_:k�������A0g�� �C���Tn[����p�Mzu $>&�Ҙ'd��"eezWGʙ���iޛv��k�L�>`A2���N�qu*�IRK~Ż{��W���� �3&���4�l-�2:5���~�7�^���|�מ3�2V�\8M~��'�(���Q�ip�%)����3X�)%<��X���Am'w�0�:�֫�b[`�+|צL���
�>�v5s���:�|�A"�&ijaS�#
q*n&O�ד[��G��U�͔*i=�����Q���� /��)̶���m�ZB���Y}�.R^���ų��S5�E�+3��Ӌ߿��uπ��^|���l���w4 }(�|}$���.�/YU�oYI����u��itȈ��tק���j�׽!�'q�ɺe�򸴊����j���a~-�M(f�p��ma�]�j�ұpsZ;e�L�d�Q�cU"�nv�eJSx�v������t9d	��w&'y�s�������¬-c�s�0|Tj\�yv��a���=��f�*4��+���Ћ�[�wn��b��8�~�=#d|��H�=�s�QA�V$z ��۟��w;k�P7$p@�FE�Vo�P��T��E�ga��G���壘ԛ�ABb/��\����/�,�������[e:�����[���C�)�c{1l�Bӂ�6Lq`�;��� т�,Ĭ�&	[�TNLX��)9S�ϩ��
�]L��h���TΔzj�5�)�%}&�#���̧��)�Y�B������"Q�����Z������}O4V��u:�mPiy"ɬ{۬�Iy�
c��1�_o��kN��N\����|F�6��cܷ�����x��h��c��%q�n�#Je
�S���ŵ�/�ֲ��)ZL	�u/��%�2����G<�ه4q�)|mr�b.��i�h�VQ���=#4OQ������f��d�)�kTֳ-q)�s����u��g���X5`�Tr>���:-�3J�/
7Q��bK-���C�ͪ�GCypGY�ROP�����ˎ��
���OIu��o+�A�#��l�UqK��ٺ�]�8[�Tٕ�hR��:siU��������W'Gv
������zd ��%�v��;B2g+�ƾ,�5�1�����]m������������u8 �5�2��!��)7}9�[��� ����hͫ�^���6�>�¡�YK\t�FS4F��[����k�Dc:�Tc�d�/��z�Y�-u��2�r��:�,k�����Ԗ�s(���,�HGc�s�{dD�n�9�CU�k�0���&/�ꉁơ˲o&4o�7���n�*|�Aḓ������6�ZY�����rrR���j@��J���$-)��r�8��S��L�AeĎk�|� E�Z�E��\��[�	�����7ͻ6�����p�'0��ï�J�ꕸ�����Hpk����w3S$-���-ࢧEʂ�CV�0��Y��u��{��0�4VG����>}�;�c�E��;�i�������+ndR�$���on�f�)����ꊬ����Z�M1o�I��5�{�=�d����a��Z"dCΐ��[�� ��4��	9���\w��7�v �#��d��zĵ,�21�YY��S�]7f�_��F#CYt��v�C�*��m�T=oM1�Z�ݦ�cv��,鱻)�1*���(�:�9}hW�%��=��	��NC=K:H�d��\���&�d�渆��1����s'BL2�FD�z·��8K�牁��L��L'yBj0�F�^�`���q���$&PYr�َ[IQj���V��h���ml���R ,����ڳ#dG�E�nq�.�E�� �c�*0E�_���(lUA�rF�C��7��RV��(� �*���f�;�?� wȞP�]c|a�}<���4��k�<_�&w{?�r�23��p0m��[�T�C��Z>P�J�t�(t����/ӀI'o���i�yQ	��?�-_�N�EI���"��[�&�=-3x-��I�{;�ꡛ��f��CNj���~�u_C ���G����w]|�P%5�m��sĻ��N��_��zT�}:������a�W���|1#�uGdǡkX��k���a#� �ctf�'�����N��xmO}2|�<ͲD�;uCLD�l	_��L*�(�mA�ٗk�0b��o�-4t̡�e�ZB�I��樼ԁ�>�yO��S=�92�ʒK�l�彞�wfV ���&;Y��1V��2v쬺]0�l�_3�u�w��ӯy�	&��Av�ul���ݧ�ܭ�Ք+���y���o�"�������]��{��5���.����s�h�v��~F����ӵ;���#�2�� $���ϱ���W�@.�G.2��b���G�3�1ǆ��7��V�d6{��DhL�s�.L�Ⱥ{Ć.U2����$kKj%�lP� �ma�O.7�*~�+���2�|��%��+q�&���;0'ݴ�h8�hOA��[I*��HCF�Sr=�_>a�D<Kv�(�xuYd��͑�٪5��8�&�h�FO�nJ���i��&��߈�ӧ'{Ś�Z}2Ë�ݗ����&O�Z��r�w������I�9Xj88��@��7�1�B�y�J�}�B],�}ȳa�Aa��>������(±�6ݚ�t�"��r"�#{z��)�����T�q�����1i{�9��Ɂ��S͌r`����>�w7�}���h��3=l2�FO3W��hea��	�3va>�Q@M��Y�I�qX	0�D>q:_(�c �|���r�M�_���M�K~�n���Zܑ���'k�IO`*Z�R�U"F�P}|>[��>���y�p�o@,8U����~�;�PeH7�!Iq3�͸������{��=@_�u1А9g���Z���T��Z^�7w��2��K���2
=�'ӷ���
�����eP)��\�؆��,�v���'��!�vlNpi)��T�%�W�glh�Dx,T�0���P���jdg�P��g�}%B3wy��@8��z�\�i�Y�%ꀦ��мdB�'��h���j�ŘsxRR���-��O���RqO�%��7�n42WSԖL�Ŋ����t|:�<�����f��[�W���Omz-�gt༕{�/���o���e����s��tp���>���a�iC������7w���0���	��ތ���a��-����Zdv����B搀�j�j N��V��ڌ����x�Բ�,���H���D�b3K:� �cD��`>�XrܐY��%�:�g��d����4��X&�E�~��Jf�b�h�=�U�e,��O�A�Dî��|��<)���-.�Nf�s�X,�/y�dJ![!�9%��1`��%O�mb*6���]�d�]�aT.�&k���>����*�kr�o�Ȱ��g���)��t4�I`c�ؘ<�NC��ۏD��LC�$)�mOR��BR������|��9e]�d!�J=����$F�R��ʶY\�����&�'OL�BuQ�K,�\1C��o���-ƕ��^F�]�n(�j��܍���ڄ��/���x>y���[D}��[ެ��>q§F��#-�$��k2S-��z�T�_�?��[K������
��Z�2!Mw\sή�������ƐY��)��k���%s!���`�]g��r��꾏�U~*�@�{�o�
�|�%z.L������yӂ?���-^UM������ӝ�K�FI��찉�+�϶��Ó�� �i@�M$%��?���0��#d?-
�'T�TbҒ�
<��'U�
UNRm�C���RۆXk��;3�oc���F����@X�]��g<љ�;�q�_yF�eV���P���N��'�(]}�1�+٣w+]C���~��HG5L��e2��3�DG���Ȥ��]��(��Hr^�N�y�Wy��	1.ǒV�N� ��	R��Q�z����U��������8����$	!d��P
N~s����Q,"�;B�bc��X��JU�p4%��Nl>>�{�=T���z��z �&H��V�Y}��8X��8�.?I|F�!5vn�7t�/�I�?�m�$O���vD�Ֆg�\er��4^p� �ktZ�R����CjS���>�,#pȏ��o5ot),�HVsؠn�O]c/��n�i��e9X�@ry���d��&���ȶ��i�n�a�W9c}s1�5L����a���{��i��V����xs�^6�'��׼��	�BI!�x��0t �����a�TE�[�ˑ���Ք=�$ ��o(봱�n���p��;�{]��[C$+����Z�O5��.���Ղ�ZbH%�y��Fr�<L�Ve(}>�r�Z�*�[�q1�����Q���dGj!v���Vmϡ���J����c�p�4�78��8�\g-7�lS����)� �����'��Un��1<��+&�<c��X.��ϕ�5����t"kT�kwg�k����u�1�}o���R�o�E�x?����$e���>���뎧��e�~^=�f2a�[+Ed�,qۃkW'�;V��*d�rbz(���I\�_�6������*O�F�0Հ2㋿���e��ݾ%P��M��G���{�|3��)�ج���d�������_��Ɂ�N�_eM�����(T�H����1J�#�,����Î�o������2U`)���y��j�. 9#�G��[e���8�5,�.���e�a5�o��L۽P�0�IQ|��W��%��P����zqV���\��D�����K��WZ�4&o9�S(�#V��jҲ���A��rɬ{tr����omބ̨�:��,凰�|��S����Ѕ����;�㉙��C�H�� ��1�jS���S���)���5�U�,���22�+~X�g568��1��p=�t�%<1�ZBhb� Rb��N@��$�b�/��!�=S{f�G���C����B�g3}��WE	��VU����>`��|�#���zD-񱮊V�w��Oi����ѶD�;��E's̥VSE�b���6d�%�y���I���N����Ck06�3�e]�c��!��g��F��R�c�ȍ�H%�~$�[�X�詍"۱�Z4�f \���n�	Ix�ʢ�_J"lMA���ְ"6���t��ɇ���({��1s���V���Y^�E^|�^�
b�OʅC<��n,����lF����}m�s`�-��	Ox&G��H���R��*�_ł�9��I��7f�ѭ6jZ�U�02�=q ��]n��q�0?^A`��9t���_E��~�������55#f��7�D�A�ǴCdR%�o���Kh(��e��W��V��~z2��fJ�y�,�$e~*+�1Ro��s�%�˜�L����LG1��-,bN_�0��c*���402�ħ?1��ƭA�Be�?�N������-�R �M�p� <�y����[@�%�]��^H0�4�������3-'%�-ܰZf�G��kL#����L6V!o~���3+�����*��+GzQ��K��b��vت	X��i��9�[�pgq�6q�a�޾C���j4�¶���Ӌ����;Ħ��:w�A�z�=G��f'9�LX���^�)�|Z];X��;)�JȰl�ު����e�CUO��g!Z���z�<�bm[Vq�>T`#A�U���N�QBmGb�w E�p.}���MX�o����K5j�>[B����2�4~sĦQuf���Ӭ�D��7ՎX	�|C��5��53�V�R�	O/�?���������s.46�#O_��H�m����ByQzԻ`�4D�����uqQvh)I��W���$�qc��E"��8U�o��}�0��Mv�]�)���2%��ˇ���L;Bx�I�(n_�-�N����;��A e��������+2O<.���U6�L��p��=�C'm>��}��6y�ӹh��Z�Pb�6�����8e���<�ӳKpCn� �!9������Klh����\#��G�>�p/����<��uw��j!x/�۳��x�.2��G$�Nw�9K��z�����5 ���gϜG?�w!K@�G�`�����5-� K�u�E�
��y�4���(�`����
���ۣ�(߸�J��g-j%I��3�ho��r��V�"�A��>P� a��w�p3.��0���Ņ��!�]ֺ��gX���H��w�������!����M��/���di�q��-i6~4���ܲ�=q��Lv�c��Ӧ�ۀ��Գz���N-.�(쉐Ÿh!�F�_��p=;�p�P�|#����03��(V�au�5�ӣFXK;���e�r��M�&&B��)<�7(��ǁER|���x��Gc��~T*FqOØ�	�_��}�y�gD�
���s*���ga���w���T��Ow:��y:���bD?i����os�K�� ��!L�2~�6���[�&�`Wg���­Z����8 Mj��3�ivC��6� �>]��ܰGW+y1�mE}��YoXO�j_�˶j���Пs����Ύ��
�k|%�>m?�8���Pu��*�]v�M�/6]�����I��W5UW^��:�wmՒ�Q�֪ڢ�6UԀ�@v���,��Viit�.W��Qsy+D��@��A��b��h�Y ������/�U7����U(���	c
xB5�00��q	%<�|čjs)��ti�D�Uݚ|���u�Z��?h}F�}�~�E�!%�+��|}�NK]�qg�� x��^u�cz4�7�+���C���ۏ�ﵘfp{	�_�$� 8nI����J��/V�������p���r*eX���-Y�I��M5��^.��5��c�eZ��6��[��`������C�%��
�K�B
�dzis�Sk���=e���nVx�{�_,#�p�,� 0<�9����'Cl��u��y2}Y����h�S���[���Þ�ٍR" �ؾ��g�m� ҃��7p;5�U��9}|LJk����-mVT͎d�����YL�m�����" :�~��y{M/1*d\(Xo$�9�x���+�,D������E��2�x��3��~�d�^���9}Hl����{@����/�M�����|�˘3N�������O��7�U�������"��mT�K�|��w�`����ؔRi*m(<��K-����H	"��u۠~�^]�J�� �sW�-�I�I²u���j>�i%ߤ��������u�tl\�m-]��S�'�/��3��7����F�1�(�;"��+cx�XJk`|P�l�,�#�2�%��q�*��S{��8$�QY���x�#ɏ/oͽ&�p�*򧕂��~�r�~R	�&t5�`�Z����w�G!,�>e�x��OY},*3��L���|ؐ5�����An09=81���_t�D%	S
�m���p�˟2���&m���T� �*�~�P�g8|Sȗ����Ӕ�Q��"�<P`��U��qfDe���I�.u�r.��1�Y�?�S����k�0F�R,�.��ۚQ[95�ޖ���cB����	�Z�;��o�xKO^<Z��e��B=+��룟*ߍ�ibB��ݱ�*�֛HKAs[�l�{H�o荽	Ï(2�=�9��A�_N\��ߗۚ�/9��	m(Ңi@�~��{A�S��s۝�v�e;Q����C(��&�~�&�-��������m�Z`�o2�
DQv�~��<�Q�*�)=��5�Yc�e��YG�mWe���#}�����鎬1bX��s�<C�z�(گֲ?��.�3î��0�P��Λ��`��X�OE�`K����_�BJk݃�
���r
���|A���x��u#�z��b9���d�'1�Ȍlҡ��y^*�ȹ�pc�(_;����b�˥�L�{�j3E������2�
�t�FÒ��W�ނB������	+�ҝ�$�ua��Wu %�lۡ�Q������cE�h�����b������W�ʇ�U��h�_p	��׭"�9��>���9W�ס oI`�g�L�V�zO��3�	���z��r�zzBd`���a8��ٺZqH������Z�7��9eī�-�n���	`)��^/I����O,��xHY2�q�Ȟ�5^�ק��B�Mn�O�GW�^c�B�O�?9�)��z�����1A�-��?�$"XP����,�w���u�1&�\����"�+I����cXN��Z�N��,ռp�1(����?mځ@�񱧈|./bA��S��YU"3!p��8؆� .����>_AƩx��G`E���j�P�fe�U����m$�F�.�O�ނ��/n�	���?�D�< 6�7�))m�v��<e���v�8�	p]zD+���K�B�0oE�ȡ��-��ķ��I; ԝ�	�ᅚ�u�>q,�9��Y{s��9C�H�}�����׸��T?v��jHw�N�lL/�-��D���o����Ո�gl�xe�P{�A�6\��<(S皭~Ҭ>#��D�ZH�B�vslwh���_��z�����Gsb�;��X���E�82Y�0?M�}i�n�	����o�%��.?h��G��ry_�G�1F˱=�b�O�2[!nxn��{��/Ϝ�:D�5�������	^"�q��D/�ꙙ<��c�l�+��dY����'{����4���8���� E^�F�%�*�Zz�h��_�m��n�W�a�����m�R�X�=�P��KZ<��Γ��`��D|���x�h�&�C��}$5ĳ�����3���W�[��J�6������.�0_�Bg�spAP^��&I�s��ڝ�*l+��s&�#����ə@�3W|�������ɖ0}dq����o����p�i)��0� �k��_�
'�p�̻�$c�9sN5�=i���˜�G� 2�&�����~�!����D��DF
9>�0����R!���NeF˕��3P,0Q"��h�q�x�{j)p��׬��ߋRg��s��¿���`�SG�'�G���;��X�2+�GY�y+6H�b���w�bV�\��&�-�5Pv$���jNfZ�i��������|Z��P�S�4�G��I��c�ށ�i�[	�T�_�����lX�W�o)���41�vג�q���n�k9t�GK�$�no�3v�[>kq+�Z��j�*�}K٩��?'z�TY[S�IB�DA��Y�:�t���(������k@�W�l}8c\ղZ��ݫ7;�I��Z�]��on�[���#f�߱�Y�����߆��V��rJ՝0��E�Y��ƽX:aP��Us����Zε�G����e�d���{��L�h֡2	YbѪB �4#I(v�9ÍMm�K-U=Ӹ�ӱ��/D�9�}@y�Zo�$r��P���łq���Ӡ���ړ�v1�F8����+���7�Uȇ�Ք���(X8O�VH�B<jA^�␁okcf�Z�����_/N���T�K��یօ�̓C�\Ѕ��e��](o���N԰�����#<{h�z�L7CUQS���A��P��Г8 �ћ�(ԍ���u�7f:X�T�h���:�X$���?Ev��fD?�ۚ!^��f�R�ܐ��2v�` gE�Ꜻ��O���#-�׭
2�ɠg�%�l�]�>�)�}4q8}�;���̲�l�X1k���d5Gk	��ΰf��s����:q9
���^V0O����;�u���r��H F21�O��3���\$�xQOO51������u�����������*ѷ�2ǹ^��s���-cu�Q�bԲ��td)o3�b2�UGUb�ĚRST`~A'�p��H�䫬��	�j,:?���s��v�܅�gd�B��r������H��
"��zɺ��m�p�n,���'7��S|�OfS�]h+=�V��*C��7�j�B�q�MhF�O����ێ52�ʰn�@��9+�n��LN��GU��a�9?���!ܒ=��DXJ�0T?q&�Vy��Wڰ�)��th(���uC��+`޳~'~[}���]�ǠA��da���g�����wj��;�\[�5 Ӂ^� -YP���-ZxM�!��Ʀ`+���?���?�F��G��D���y)��7�K����*4F���'�ҧ���a���{xF������P�[.��0U�*LX���.4��;�_(2�GkA!�N�#��%{���duT�36dtF�XK.�4�Q���o�I6�z�p9J��I@�	����=NV����X��8�$�:,���E�mN|洣�j<�u"1ֲ�����{ϴ�bT@���]��Ƅ��̄5��3�Y��O� ��R����t��f���R�zK\����.7�"���OlK�d� �ܦӹ�&&?.�]Q�'%,�Ar�b�6 �&F���a�)#�S��\l|!!B�$4� �*ܙ!e�z�No,�V윴����O��(��	em�� �a�Jd*t[6��K��f|���DpJ$���&��r���"��b���$89`�J0�����(���n �5n�6�Q��A@m��X���R�dKHI�?3���Jݢn������8_��AU�K���t��d�}������C��[������J���@��}�eZ�'0�P��.��ݴ���!:u\�9Y͵u�H�j*P�Kc���ǼȠL��n������5���s֙[9����WR�O����m������_E12��k��T�ð�fD�C�����01:��m'�T�@9I�3<\\wH��(!A��XY����#���P�����'�W(g�
�_�cBJ����/�Q>d!�?�Q9n��fC��K�t���mt���cղht��$�a� ���諗��5�S��7M?��%$g^A��w�8w���y��_���4�O�|֩�2����o��*D�?�8����ؔ���i|r#1ZQ�h%�&����]�^��E��5��(˝Q4��Ho�$�!)��I��S���O�����^�`PD��.x鿵��e_Ayq�˿�4$���(��U0����|x���6O�ZB���]���u���9�,�rOE����%�����{�
Yqυv�@��R��B�<�A�E�8�����L1.��[<�h����;����Tp�j&�=Y���3�_g����.�\l���n��!c�M�K^J&"#:̑�!�YN�)�hM5���8��c�Hz��Ϧ��z�� ����r;���kz��a͌j��f�v�? �WYU������,Uv�S��z�{
����j�Z6���FZo�Ͱ���q���}p&��TQ��$xi�F��w=ƛ�Hᆉ/o�:��fڲy��C{���!J-E���g�)S����GSv�m�2oz�6��r�pXZT�׼>��B�9�M�H�\0��ev�/��vʁ�h  ���h�ߏ1Yp;ٻo	)g��1�6$�P�C��B�]���G�����]3��h<,&%#Cdxۙ��v���=G]���H&"VBIhp��;t��͒�q~�o��`�v��{�Rj��Y9���	e$ѥ��FԚϵR��ڞr�	�`9�L��������hv-�%������������Nn�C�6���TG��"N;wq)��z�t Pbx�6Jy��v���6+���ox�s4�+v�$o����x�=�ajI���_&�/���+���b/��L�����7�z�������J�G(�Mt��2f��U�i�h\9A�틤�V��me����M��Kb���+��['*pP��|�EZt��n�zM�����hW��J:�K��3�V-�)�1�O���jS�5;��Z�u��S�"UZJr>��}��w增��K%�o"��=D��7�♷P�k������P5��!M(�5w<���#=�
���آ�
���;�>�l�O�����G)�TC�=�C��Ϧ��;,�����I_�XP�ZuL�AR�����kGͥj�(�_��	:�eTD�;���S�+b�/c��lq��N$�R}]:͘O��z��4�M��6^W.�j����;���	�-�o?n3X������v�ɻb�������Vy�"�1�R�{STS�*t�~'@�'0�#�R�Oh�p5G�gΗ	��nNS�zoV�^/R�E�	�,1X�5���2v!���t�̠!5f����X�i�/��#R�9a֬��3[��!)�����Y��i�ңGUx�G�s���/<_1��;�q���B3�jv3FZ�?N�t�g���1��?'I+F��*���R�Ś`S>��k8�B���#C���l���AM:��*��s	x�'�)��]��f��@�,�Q�N�j��PR��֠㠗X
i����H�����Q��2[���:zyBNC޲�q������l������YHX2ů�Qp*�(a�K9C��K�E�ݚ�R;�Z7X��?�N��v��O���%�Aų��z�i��0�ʞ��	����R�-�R�����P4��n�#���F���Xp�]�<�>j��fH^�:�� b'�qouD"�)�`ǚ��
�N��O&��/Ҍ�=�3�GX!��Y�`��C�lk�%<��r\d|�!}�ql�ER�ho���;$�Ё���Rʯ��~r	b{�ZPH���@�+���c,}6h���u*q��!�aR,L�\��zP1&��c�H�;�(%�6�}��WjQ_����������7Va����xV4�󌍳#	V��Tj�g�6@��sEٱ�w�,<�E���g��u��Vp��i���S��
��LɆ����8­�i��՗���y��+�V�[!NB��mhܣCѸ��X� �`�(&�������C�e����ى��Kw�Ÿ)��+c���6���H�	�Z��\@L�H\'���7�{�IN}j���9C�Zo�X$�� ƕ,Op�4�a�ء���вf�TU���)��י9ZR" ����s����V˒Ȃy�&#��|2PH�~aκ�u��o�|�ܱ�!^�s�����pTzFu��A�IZ��N���g�X��V|{�+C���L���`I���y�h����W��X�DG�W��e}�0�O�t8Ƌ��\Bf�4�0�?��+��*üKW���Q�Q$$NI�˸p�"�'q q;�+ƹ�P��õ\���{ш��5��
�$�1�<�U�~�d
���M���� ����,��'�fl����]>M�͆r�K�~���e��עK��zJX���ǵ~�{}Ⱦ$�y�������"����uJ�1ڭ)��q��lA��˹i"��=���!V��?�H���Wۓ�����ԁ_��L
~���P3,wt�r�σ�]�C��>*�;Fw�@펍���SB�x��on�l��e����f�;J13j���{���T=�ݣ�h[AϥyqW's� ��vp�e��-�9a������̤gOv�����2�g&����u^�e� ���C-�
��)wT���F���t�j�viU���Y�0�c/;����~�4HT%�6���p�I���Mp��	�]h�&%�F�D�)�W�[��7uũ�+Q]1�DuL!5
m{s=��4qtȿ�|5�-f@y�ݱ$gݚ��U��K��s�E(�͖S��q�3�+Úe���"�d�̿����!"�:m��J��U	���
帮D��0�`5'#�i$f�5/�`U^^��'s�*l��}q�huJXR��d�GЧCH��>.��j�L�A�� I�(��{خ��*2`��*�/��f���[���^��C-�2�s������8��Vh���(�Un���N�U��*P��f�%��m���Z5&���J��/1�����4���䄫�:���7���Q���'���2L�M�{]t�٬���C:�&9�KJK�u�DG��R�vW���\H�����R�8E����$��\��Mr�"��1�SU�W:��Q8�/b���=2����l���KD:La�������ԢU�a��l2e�bU	h$�a���d�a�L���xi^��G%�PX,�W�0�e1S�tF8����@��6��@b=��BT����V���G'��GMJf������qs�ݓ0�y/���K���tqWDAs�?���F���;��'��e���gv�[U�6� �Е��9�Gd�Q�xA����L�����^�zh�vy:'gO��wk{p7���nlB%t@ܽ��N��ЮJ�h��I^�Z1���ȡx>41�ᵜ�G,=�u�6ν��H��@GᅴT�����Sٹ�;{��p:#��ƈf��F|��R�y^�&W�����e�Ca�>o���ۑɋ�.7�I䫏�� Ĭ?�ƈ�Ҍ�	�@5B�2)|@C���o�>݁u<	��Xʵ��`-QAo�(r�'�*�6��ׁ�d%}l�?%�$BLl�[�
��|EI�H��t��u�=	��Xy`��İ{	O���;�T��H6�ﳥ�a�rk��t,�����1Z���_~��<�UF��n6E]|�(�����z"�C܉����
O����	.g�=���"���E�Բ<�1�r3�x`�~�+�(��Nm8
��$�M��jD����7wv�J��ö%����dK;ӓ]0��/�Jb�"˧�F
s[]�����2��U�/;��4��t�<j�P�tMM�������L��ԫ@h����~Q%��U�W@����>}hi��}U��V!��\&,��(�N�u�c`AH�Ƀ�fv��-[���Eevԣ#�O��}�$�4�s�P7��E�sNb���\.I޴s��S�D����q=^"����"�^�7���V�z�kEO�.�*-�K{������`�?�<Y���2���j[���	��W��j}�!�W;�5W����$ae{�L�5�j��9������I�]�.n�#(����� �����j_��������u晿PߠAP��6���(_����
`?��
u�y�*S�����5�
����"�NU���vs�_�z���m �qp�VÊO0P��EEg�(�Y�^�]U��y;�6��֋5�۴�w����pH��6t�~�_?/C�w�>J�~-�Nq���+x���1e�?�]��7���L��0@c/=��]!~nVW\���l�Bg�T��&CCg^��I�s��'�t��$��1�Z����;_VGS�X��$e��+%J%�kG� �BR<���x��Rn4��u�YE�+�|i�GI�B?�]��X՘H¤����h� fы�jkC��c���~hqw�q?�Mu���Yqf'J���@=:l���%��.%������i�h �VH:��/vА�fWj�ë��縵[���Z���Ѝ-���{T�� w�`J?� _}w׉� u������~K��y ��qN�����f����^���i�Y���g��
d89H_�?)�/}^V�F���J���dv�Cq�������w�˔kH��B��h��S:VRH(�ο��ϓ�0�id+�1D�fP�hs��f��ږt��d 艱�������輈��zlwz;*�~%�\�L��q��@#^�6U�7 f0{���֭�nf��o(=��.m&� Z�A��U袶"ƻ��>��[c�8��ru-��B��ӳ��Wf��7F�D�y豿2H`1��Os9���8)=#�V����5�y�sV!NEfzt�d�7���w$�BЩX��+
]���N5;����Ai����ڴ\���×��5�ga�OW��n�E�jvWU�i��e&p[C��q�DγYd0����h�IY�PgK�*��z�7F���UV�)��0�%��T���@�(^�u��� A�QJ׎ء|���NL욨�Z�ӷc�Ą$^�}�g�*ͨ�P�����0	�A�ƃ�^'���9�
.��圀�{�O�5��QH���D�K�v;Db�Z�k��TQ����X:EH�!F�U�t,��O�_��
~2u}�	���7���B�+�I��Hq��,��m"˻�N)�`�\
��2��DM*"6[�!�|�L(��Z��O��>湝��_h9�wF�v��p�G�H1s�����I�0^�2����t��{*{ 9,b���E��צ�Ƀ�la�k�}����N�Pb��\������|&��G>��8acE������]L�� ��z@��&뽺�7�j�IQ�P/�M���Sv� r��܌U���1�1�Y
��:��n�`�̋6�7AR��OX)���ISH�@&�q��	M�M�^㑎e��=�M.�&��u�@�I�^1'$�E�/u��P.�Ǚ/��։��E���1��&�Q��p��-'V�E�0��kS�g�k�ZtSs��]���X��16���rt�5�3���<��!�;����')�n�(�`��d�yc��������h'���WzI*�s	���z��g���#O���@Jo���s���&��J�E�_+��f��T��a�e��[S.�E���k�t`�v�p� �Y����?\q9�:*{=��
�|-t^T�R�۾"3oNH`Gn�u�s:ݦ���ʿGf ��ѷ�y6������x$~��6����+ܷ���Co�w��ש�WJM$�i�Q��\�c����9k�;���(k�C�$�w�`�+�U9؇s1i���a�|Rha������b��1��9D�Ԁ�}�����XhƐH��:��<MU	�X���Vd�o" G�B�[����	���T�%��Dw��A���t\3��Mf=�y3�%@�������x�w�(Y��}4O�D���=��[f�D1ص�i"�C	\��j��bY��1�,������r,��y;v�1�����@�̈f�wO����Y�m��,���� �tߗ�	�%$���QɃ��U�H�cc,�#���}<|/	"�pof������0��g��۷��Ƞy��h���j9�־�ք���ȣ��ys����񪄒�SR��� �Ş�Ӑ~C�R@����F����a�0����7M�Iq���xC!����(��<�d>�?�9�+@0��	����-�6���<+Oe�^��&��ڂ�E�B��B*?�uG������c�I�+W����3T*jQ��Aӻ�'������ݚk�};�I"��^+���L\*C�7�H�ox��?
T�nw�g���b9Ij��H����Sv���K����ӭ��'��eD����Ӣ��r��"]������k�,����Gx��$j�Dz{��ɳ�$B�T'(NX׽���Q�,���9����@�~p
1}J����&| �D�{�a�
���X�F�E,�m���۷0���	������S�dJ��O1n��69�d&���Nۑb��f�.g����
��U^��қi��6>�!��'�~�PW��L��)qAm�P� pM�h�2+���>�K�1���-�0��೘ 1�f�k#x+�U���y�W�7V���|�Gs��Փ=�gO�3���$�®*,�o�i�����-|����_K�=�u}Z��#�����	�H�!�fR5;!���l��S�ƸXG�3�@��Ϻ�Д_��7G�Z��ڑ9*\��� {)&�"��;��p��谁&g֢X�a�3��E�����#�t��r!���o�i���|����4w��&t����y�r�Tu(�g����â;���"b,}�E�
�Y`'*�����Md�q��k�} ��L�û�G���a�
���V� �ij�z�.����~�K-���Q��ee4�z��3iŨ���!�K1�+m��,�BH�x0���dE�T+�9���Qw*F���巈����
��d>�T0�C� {�W�/�gC�_��-�f2-�2ɫT��~�
���
��Y�U@j�W�,��ޮ�]�����X5Hن�x��J!���x�%V���0q�-���F��p�R��H�l IQ���-ED˲��pa��p�!v�M�g��a��E�@��x����9&bE�z����1VHE�ݚ��j��k,-ߖ��_�{�����*PJ��ݒ����+��,�9��V��NT��_6<���jS��KOK=ىD�h�.��K��������'H�\�!}�Rj�n����̆�
	��^����'c���^�눊�(�6�=f�f�(]k��jF����O�򇼣������wsA]��hǜ��t����Gи��sG$u�j�T����&f�~�ŞHd��pLw���WM�Y�	F�1@(\�l<�� u�/�T���9/��`����_ؓ˞D.����k]�jA^�
:�+ǑF\��+˯�� 7n�
2O7�� �T��jtk=.�a|�Er�[pk�&�ȅ�]�����A/����Z�F�G�-|[��9�d+ݼ�gB�ay���d��J�RG�>�c
6��,���p1��#��^��9��L�{}���|�N�t��K0�݅}MZ���C�f��	8rzo�1��(�����%]���=ĝ�s���񔤀���j�n|�c��ش�Jq������1>��q#WA=PN��ּ�	I�jfs����m��o�l�<�iP2WB9' *	8q�S{��)}�4� ��@��v �5[ATD��R,aO�b�%���0@0���|TТ�3�����~�e�����g�N�LY�����Ih�{C�Zr"ϑE��5�^�?�Q�2!���c:v�}��z��k3" �<�4��i��.tǺ6�FD��R��o�~����q==2��S�i�r�J�݁A�}/�i�Й�LhY��������1^,�cW��Ɣ������i�-<pPHu� �Z�ʄ�o��zN��k���ƾ�]jIO�u|�WbW��KvSbZ([47G��?r�}NM��^��'btz�62��7�'6A�k���Jo>k^�*������Q�VT���A�(�?��{��<�����+?�w-}�������CO$�FՍ�1���w�\Tn/3W*��Qp�
7�D�,�ۥ+.�Ҭ��s��I�)���z�[�]�T�L)m;�~�\交�m]���L��ڶ(?ğ/�Dgt�Ʃ�9���%��'ZA�jb�b$����ʀ}<̟8+��n�~�0,-�:��h��X�cXOޱ��%�}1�e�x�a�{�����Дᙩ\mJ]�F�ǎ��F.��:đ[zb��a��,Y)��6�=���\4������.���6����W�F�FSHX�T
��n<秇єy��A�ƻ��S�y��&�i$"���f�;
N��`|��M��0ǝ�J-���ǩ})8��{X�o��KK�����B_�ĸq����U�G�B�1������� D�-?Y������BH�Z�bS�W�f"�>�Ό,^�e����R��k��6�\�\�+�eL�"�5���f#{���"�ϯ�Ѡ��*�-���X-n�bYf�jt��o�eb)�ۅ:����G�S�Y���S8��@��ѐ9^����c�'��m:�DnVsb��<?��U���g�r�>y�Scs�XՅ�ŚQ���>J�U��.c�Uܨ_�%��ZU0����:����&h����Nl�S��BP�U �b�=��.F�+R{](����t"��f��(��Tn=�%ՅUoO4Dr��H;���p;A|\z�2ndb�pNW
�Iqf������<�\��)=~СVg`:�bԂ�)�"��- �i��RܦL[Z�0�q��ɲ�R5��f>PAe�^_�&i�bx����ӡ'��$�:;ZSx-i~�j��&έ��v�Vf�{;O�㟭NG'��:u1|g�d-ݪ;\���܂��Ja饺vСFBp�Z�'ǃ�ΧqѶ�-��(~��9L�8W�u�$6Z,������"�,��޾��>@��4ܰ�	,���tt�v� ���y\���Ԃ�:9�~��s�V�xN��
?5"��BhF(�~(!]��&Xu��w�Du![�]*X�i#u5y���ؑDVr�5.7S�ƹ��r<f�\M�:+�r8�50��J�%=z2�G<ŷUk]��
��0l�������~*���8��r%�S�s��r %Z,�M�ˌ��oR���Ae�`���8��d��5�,5Cu���o�u����I�F��2�˩7�7s�"�?�LB/@*T,�ĸ�$^l�M���w�-�����O�L���U\b^�aa:�IPVq��z�Ϥ�`��ߩ��bhؙ#���u�'7���MV�\ݙ�7be�S"�������삞���������a���8bW��إ���>��c�j����r:(DY`e�K�7=D��$�(�4�"4�D��h�►d��'�Ry�1P;��O�����)~:�L���NX����l򾲓H�Q��J��石�̈́n�@T5���.}hx.��;8�-�#�OS��,d����X[���#H`����v��}�Q�i�(�3�F���������۹�B����qEy6��<�
S<��|��u5�1akwCBe��@�,~m�w�6���葱�O���G)��Ւ��؄%�{m�m����7�r��+�*�7���^~�K3��!���ɏa�G�i��� �����Xy�孛��^C2����'WP��sܺ�'<,SE����v0�D��r�����A�<��e�����3��5���߸���8�s�?.�O�ǭ�a ��"�������H|��f�j��Ɯ��E���QHH+��Q���gI��su��U�C%���&��t��+�͚:t��34ֆ�?�"�� Ս�xJ���T3����p`m�<���'Dnր������4�O�8ـ0�xX�c�*�������:x �^���Ө��jQc�cz����-��?�h*��,��}KtB��+�7ij=>�K���
�P�옰��\�;�n�?�`~�6���Fh��a����D�`d�^a/3�$�\*���+�	��?c1����h���YJ��t�p��9�փ|�&j�"%�M��0�(b<aH[��C���9<Vc�bw�H��o�S�˿1L�x�?�x����M���Jr���*rSOJB2��N���ڊl鿟1�?��Ym��J��o��g?��hȁd[b+1�(��.ym̚����7;5�_-O��2��@07A���J����Nj�e��C2��!Kqǣ�+�2H&q�Yb�J+��.)"��nԢ9F1t��K��ow����U�ӛ��(2�4��%���_Hq[4����lZ�2u���/]� f�[��+auB���b�Z�|���/a[PՆ�T� ���[���p64�d\�Qd�/@��3@� I����3��L�9#s�o�:ܡbZ��c��'S ��^@"u#H��;;���u/��{�a.-� ��D�h;)NƬ���k�ۀ�ڢ���5���Ŝ�\����Z�=�^���$Uw��~���ٮ1�!L��;n���u�1���G�(H5O�Uxo�Ρ\]�����{�M��視�[����$w�u΃�B#��:В�}�yD��Lk�]e���p��w���gJ��}:5l�@ߙx�.o�:����C�+1�v��a��3��[b�Yuo;��Z!$w�'�P���%$���Y�A���=Op���(_���5ds� �H��Le0��}�V�h�Z�&�Jk��C~5�򪭛?�K|�����ϋ�̯Z#���H��͑�7�~��=�ٛ7.@J�4��"��3Vk���Be^u*��Z�0S�R'g�=,f�HR��R6a�Ũ�^�F��3v��B}�= `$ъ!�i�ǲ����+J�g�q�)z��>�Qe׶��}����Ys#Q��_�J�?�QՌ������ѿJ�9���?矞L<JR����	8n����T�b�3xoHEJ��Z����0�öT,Ii�^��R�� �6C��V%��T¤�]����#��ώ�#��i�~5Z,����KzS*C��::֏����1p
L=����T/o΁{H� ��\��ʨsի�}��fC>��N��i��O5�ʕ���$e:	FWJ�N��k ���߹𦐥�9D_ޡ]2Ԧ�K[v�&�Tl*�������lWs��8Av�O��P��XO�D���v�G@g)�e3\|�ʦ\wƁ��=�6�2qNPgljl���ҕ1�N�_�=���[��=�̖Ď`�`�ia&c��e�ܝ� �Vm-a���S�`���q��3�E����tcpv�`I�8�ooS`�15dp�ϮR���~E#@������=R'.�۶b\�>�FN��J�T�i�i�b�?Ǣ��U/),�)V�3��{�6���)�j�L��z�i6���!D~ѩz�Z6�V݃���=[���B+'%B�f;D���!M<]�M/�N*k�=A.����ղ�k�	�����ϽQx\"4dql�:0���1�/oRh����a�'�4`�\�h��X��p���@v���3J��Ѳ����E���X��*8_�h��:6b9��.ueIY;�Gv�j�<?����>
�թ�B�!�^6�A�u�;m�S�'U��F�զ���E�G�(F��=�Q!���ո�mw���[���!���!]"�V�Ziz�~�:��Π5PT}<��"x ��6y
��
0O*�Vw2�̜�>3J�N.F꧹�2�,=C:���6���v�>p�{�诟��˫�	� i=�[0�EnN�鞯������j�:`��W/�@0!j=��c�����YA�Z�p�M �f�\�=��E=&:uqK<��jo��	�P�RyRi���1��f��"z�%�2P�(��dhBd�RNlvw�w����	b���&��w�2�6-��w_<���g��ԂtZa��/���^1`�PAf5�޺z )|����a4`/�o���5Ң��{�`7�(f��7p���%s��V���=�|kI�5f!Z�#�q)�"�cgj@�:f�<�=�3�F-n�d�S2KŒ�9�N����M'eݾ�x�M������XF�����-��X�) ��>_y���
I�`�4z7ڝ���O��A��%���J���p7��]�--J��Ջ��xF�
�������^*c�a�9{��Ci;�c���H2_������wY�Uz�����Z���a��I�����M@J{��J��0OjZ�@�~�����R���7�3O������H����5�C�ea�wS��bWIB�F;۬_�;j6�F�7�Dt��1{��{�^I�����5�1���-A���3TZUT��n���)�3���O�[�?[����h3����n����P�w֥ރlyD�^����c³�Lڋ|K���<D3��;J����~���ZR����$~���H�f�i2�M��$�sWс��]���r��ҊOSh����2�R��Y�"#[�:��y��[.�A��bx�XƘ���[��Ќ�d�B�Md��s�m1�ڣ/�y�ﮎ��FO�^��V���F��y��/������?9�y���#t�j��A�H�QP�7���t�cjS?n����X���*�OEߧ��A��{��	�ڝ�-�6ɘ�;��Wy�����}ڱ֧����w�l��j�I�{L!-IY������K��B�V�o���T�t�����=}�5�aӲ�rk�	���7骁̓�{0�'������v����?�"�fϠBgHǔ��׀MJ9D�NѺl?~d��:��'�`a9�̞cO�}i�>i���w)�O���j�9�3�C���&6����������c� ~y��� ����f蛫��3o��g6�6�D�g^t[���������5�)�JGk�O�4�Oh�ņo��!��B��{����hu�C-p<��(`y�gid�-y�RE���{42J��M-�c��%N���8>|R� �~�	���80�I���L�*��eqkyIn%��vw�X�ѭZ�:�Hz�ѡp�-v[� |8�If�Ϩ1�K���p��hQ�pZt�<l�u��#���+�ڝ��i1����
wYr_.��
�U�u��m����5A��<yOr=IȘ@<?�k���f+PC�sU�s�K�w��,�p\�QF����c���G�b �E�%��3�(����6���:�_�gP$�U���[�'W�'3o
=�D�	0�W�j;��6Qeg{� �w�b�i�t�%�Ǉ��4#����֜K�"ߑr3�y�[�C޾�w/�׽a\s><w�`%ȉ{��"�����y1ayl,�Q�^�j�0X�H:]��N���~l���E�6��y��;W���bߨ0*����+���V�V{'_o�K��l���_bP���'�x����f�CXՍ[�Z�L{�^�C���%g��A����}���?L�۝%rl�5,,�|tx¹!���Z�&�a�
��y|�ٌ���xVW&(�Qj���m��b�?){+���^�A��t�؆H+7>d��B�.6�G�kH��������)�:I5%v̉��:Ѝ�qIcI)���[뱦�)ϧO�*���X8��-��$��O��™���/�e�%1>����S��� �.�bf���w�SFf����y�����W	��FG�m�p<ci�n4RSԬ7�h�����u�,���d�t�� j,�n}���J�*�FnlT��uw!t�8�����m�X���O�	�[ժ=?~#�lA�K7,�f��[�E�w����U�2˨�|=Z�����*���@h�]���֔�j��TR�s�U�8��8��;���� J��+r����
�o�kX� X-(=�C/*�3/�F� ��C-�2dx����K�>!��Ʌ�6֡��	�M�CW�6��"y��ӌd��g�]z�s?����E��ę�����45��������F���p�`A1�4�ws��C"ʴ��&��@ue�.F�Ξ�`@���}�b4o��n��&��<��wb�񾁖5���(X'�P�otj�#Z�J�IC���BU|��w�(uuS���n��bh��&=w�o<N�J��O���n�{��~�܋HV-��D�d�z�z�嵎�p�� �;�Ի�������=��^g�@2f�������EjΟ'21��8�w2��Yq��!�äF��j���\��=p�)�H)���D��9ڡ��-�G��;1:2�Ҧ�k�CI?��"����e-�^�w%��[b��������U��z$�@�_{ )vџ���Q�)4�R�DG����{���zF�L���d���{�~2{)���'�G6�u����FAĜ���_mjC���l��EO�`Q>$te�����գM	���Gf�'����x���m<��u)FK��O���8�AN��]�ꆇE$����;_GK��
{���*c�:�2����e��ƹ��Y�z=���a�4;;�^X��g�h8J���M�v��#埁��tG�?�ɛ�1�6�*̾@7�<����Pn U�efmEs�x:��~�拫,�����D�<��C�z��}��Um�ϴ�+'},:ȍ�E�\9P���ȕ;�=X���H�̇UH �*+��!LS>��Y�b�3��h���l���;��G;�O���c.��:�cŌ��.�<{_F߈���:�B���s����F��2�W��8�gi����G�Ǚ/�d�	����I"�&+���w��M�B�j�/{�h1���Za��%:U�77PO�1���z7T�O�pd�����z�k�G�kH���#���
����^�A��rк���a�Cݷ�<;�e�׫Ǚ�j��,Q(Q��p���G��~�nt�U6ԍS�2s�����tQcBQp�����dr!����2:�M*ߞp��%����O�����m5���pj�hq0h��
�9_�ڥu�3U���s����'�'_]�dB�>�&�Y�D�k�ч��ٯs�g��5��A���O��los`�@9����XOKU�~q�>
dIj�w��s�0���\`����G!��/\�;=<� ��;��?�
3IԬ:�n>���)��� P{��UiiE��SD��j�!s��U�ԗ_�r��"z��A�oV(ҹ����KLL|���G_��fd��.B��,Xp0rz��"��T������~?����<�yʢW}f�� 0?�8^��<�w�%Y�H,k&���q'�Z�]����%4�P�X���]�2�V~i�lv{ �{C���O��N�P)T�L��~��W������H@� �����I�?E�I�)�o�W}d,�m�tõ/V{�.'ifg:^Y[�n��F܎�?9JDQr���ȉ���i���bY�iW�'��Z�7M�a��Tf��ˈb'���5#A{ηA'M�HnE�����a��A>��8��v���yLWY� ����ż�&��s�����=.�djJ�
-��yn�~�b�Yr��QZ� ��(��ͥ������=����z=��[�73��Z�&�C��'�u�������`Pf���[v����I��W���ز�/`m ��柳�G����&�G=��a��,c�2M=q.0�*a�$��s�tvpb�9M�z6xe?�Gc:���S�D�~|��?)�k��Y�"�*�/�Gꍄ�������'�X��Yk+�WE6���+�2z>4qY���r�_�Xf���p�v��O���㺆:�!��x�P�����[�RgF�49��<R�D>.�<նM����ڌPwё.�q���Ԃs�  �"u�^��x7�t&�ŗV9t�?ꖼ<��#K�UZ�L�k��k"{��'��H����ށT���H�})��J+z�/��rH�N�[��G�崻f<��8s.(Zj�B�z�*��n��:Hm-a��.�W�C���c��d�^�m�̏fg;������y.`�'���J�%o�xX.�^��P2�\:1��Iq r�DrJ6���Yv �.
����"��N��mf�g����^̽O3O���P(�xW��=%S=ԅ��Yfs�������ح��{8�Վ/9i������`��|��LG�?��g �F���w\�F ��qfl����[ZN�&Z�Slʳ�V ���[��P$b�����u%s��{A�<9l�&�K�i7�)�1^��H�"��qNM�k��5�CwJ��B�*�xM1p�C�s瀜>�2�F:5�z;/Q�[�w�G7/�/�?�F�_�,���e#�-|�'��e�6�3#C�~/f	z#�P��!qah��`�L��M}�����?�w� V�潎�`e����Om�﵃�c\�K��<]� ;;�S��p���;��5��ݓ��.�l;��&����tҐ	��`���C0J;���<�Q�/�����z-�!�g �4��"�CFB����������;��E6@�0�#���F"�C���h>�d�$���W`b���E|uG�p@:����r���Azece�³|i���͆���[Ҩ�]L�J��BvFo^�K�ϕܺy�gHg ���0:�$^���0�0�ve��P�5��2�������y���'>�է���k���:{��B\�Q���N/몾�1�O.���1���S������ر�Ȍc��H� 
	�DF�Ou�����P��^~��ØU�y����fR�T��U�Kc+~���h!��x-��l��T�I�O�އ7|։�8܆]��z��ͼ�ލ�/�u���?��~H҉�d�\�J����}B��k�Q.e<�P;�4�<l��,��.��$�7���	��nJ�pM��K�������+#�w��f�,Ar\��4�߁��G��R������A�5a��
�O�D�붍���,'9�r�i�G쥤٩=�C��h� ��Z&���V�SJ��rW^V�JK�G���~�����0��'���D0��k��%�&�?�8l�4��^�;��)�� ���K�ޏ������pt���h�7qZ���:^��z�uLiA�7�y>��u��,F=�3�'$��5)&N]�����)��G�?��(��o�V��Qƚ$��3���ьM�pv��pF^����:�b)��� �|���v8u��!�|��P�Y/C��q�*cM�V�V�
62�2�p�rx���� H%&A�-�����2>�lxz9�e��W��J˂��/Ks�O}�eb��z���+��4�����S#�Ӈ}�-k�V���܀�H*O��Q�Cז�0�"�h����vg((�>E[<`��$��Ļb���e�?@KX9Dho=����kS�O\���k��3!���
��@k�^�13L��M��s��a�t�p�Q�fێ��i�
]�a맊��=4i}P#x�[(�Ryu��VԡR'P�FR�5��ʠdg�7�c���aʥfF�'F'h�B���?���q�ʭ�GS]ΐ$���������wQ�ܛ�:�z�C��� j�6�P?0�bY/x�jV��Q;�6o0�!IjV�4mv��y�*R�a����~�9$Ι?�cG:41�۔!��ަf���� Y8xV޾� ��K~��/�m?>`=Z� -+h���o<rb���ǅ��
W����m��W4����v�L�8�֟�on���C�xV���6�9�G(v=n��Q9��9��R�
Ŵ�a�q�J��nǑ�Y�	�1e�kk<�׻8�|�V,�@S�M�)\�
C"����h9M]�-v ��=}�`��-p�E��==t�J���)�\Ռ.�3��	�Ԅ�.�ö����o���1c���NZ޵��573ٿ}s�����t���M.��M���~�?�7\Q��_����`n���8c�%��.Y�	��D|+�7+�]���'�	�6/42\{(dk��?�m��%���2CR��3<�BDwg>5���!�#N�bn-�l�5�ێ���٠�=0ﰡ��̗~��Y��%����h��ty�C�J��.�k��҇s�����	��c���ɷ���O��4�j��P(Ds����rk��%�x�l���c���v�N!�ے�&|�S���Go������Kr��e8G^K�X��)��P4�VC�Ą;�y*g�[%axهW9J>GJH�]�mJ�i|�<���u~O|N<2�gf&�ʉ���w���lR�B����?@�PX��,f�b�#���p���W�.�Q��`�u��d��/�L�ABN;�m����`�<H>���a�nnH�� Dlqt�.Ap�vE�����d!>���_Փ�1�Z�i;��4˗v��=��t�,x�X�%�Vlb�e���E�p0;��=R�0cI�O@>	���"8ѮŜ��zہ��`s�����A�"�Z�J�3/Ӭ�"X@������S�G�`���5l`�Kf����iW��v{i\�z�F��P�����o8��0*?��2Om5Pc�#.2wJ뿲��F���m� �n����:� �0]���0�gTi]�0QX0�A�nԩ��?�$p:���H��=8B��)���l�����<�4r �u����O�/2^-\d�?�m��<=�%��T�U�o��'YV��4q���9V��U��h����q}�*���(*/����$�{3�����X��J�b�?e��QN��`l��Ta��[Bn�J�mP�Q����#'��k�$���,�Z�Pi BB,��Th$1l�ۖ�U��7ӓ(qu0����p�љ�����s����[�� ����q(<�Q��L7{��a�$5]�otM��0+��i�v���7X��:o��@ñ����47=�x���g;���$�L��~O}�Ί��w��nT�MQ<�����2���t�UQL�I5l!�k_�z��`�\8�j��V�H�?|%ߗ����>#JXh���m�tw�sCe�b�F�t���c0�Q��-�a<쇩����d+�e]W9@y��Z\�ܾ�J>b���N%5�����VF��f�q���+�22@<^����m�>�x�vDj��	|>�0l�Y��֋�_���I�	����G��\q��^=a��88��L�����5:��L���6�3Ik��rv9B��� =sJb���vYm�;��-��:
G*#�\g�E~�~=]��X��������o�t.���'f�湌�$���T¯��j��3��4A&Ӛ3��E�����`�Qrz��2p��4�R�*D����G� h}z#��s�G^�a0 ����*�@�\گ"��nQ��7`����(��J��V��*�p�B='�E2=�S>���V���珪 ˂�R�1n�o��{�Y4��ظbyl0x�ءI�*3eKW'�BJ�>��Uy��5(`�0�	w�J�u�^�d�*�^���	M��;�i�k�n�c�����#~�k@u��B.ҕ�Ht�k=M��ϙPA{�����CMS��2���\�cBF$tߎ��e�0ǊOL���Fcm�$d?c�lW�f�c<����L��q���(�}W:~����Y`,��>41�OJ��^ �2�t�^t���Z��vg=��,B\Լ����'DS�7���ze�b�d�(s逐d�;l��Օ���q��nA�\�j g��P��/A|~�^��Q��w���_|���C�o�-@J:�.�R�K���#����ܧ��<Cc�M@c�$ �m/�bUT:Ml�<�U+��Q7����tc����p\�����ux�[���f*R��VR�
N�["'Ƞ~��`�L��	h�M
��T}�4g���;�-�~y�^נtx�Tk/Kl���U�S�iC�9=��Í�7�}C���%\JL;����-&�6"�K�Z�A��ϯ���Ӷj�9���	�X)�z�XA P.?'ԉ��Ȱ��H� ����Ͼ c����yNn������}^$Տ[���(��&���V�P��[3����-�����~Q����=�#-�����E��-��s\�P�u�q�y�C��#)e�7`���R͹�~h'�Z�:�����0��r�����$�/��E,F�R�������7�Y�@й���0%v�ɴi���D�+���I���i:v@�C%�����U�An.ޠ�y(4�{�q%���7q"��\�\ۑ8YZݙ���=I�CfC.�T Ha~z�S�EF��w]��Zl[��g��g� �^��R �v��.�,<͠��tt!P�z��`Cx���f�X�"Lv0ddk���(�Y}�˵R��!�Xo�����i�ɞ��s���d7N<�~�y�m ����N�<h.�e�P�[4 ���#�C��(�J�r@��ph0e@*!?��|F˿:�\�{q7Rd�t| #w���_G�E��Z��2�7ˈ�p�{���'f�)�BѓXp���.�JC�S��1�� ��_�C���p�����莱UG��9�q�ݑ�y�s��+�yN[��i�f����]�w�#^�4c�s�*~�Hƙ�SO�=Cy.�.�]�C�C����p G�U�h�+b�Ρ��8�o��+�ٕ�p�Y?	�s<�<w��G��Ƿ�J���4���%! �_Ȍ����l�Jr�����	�4�[�����n�I\%X
�K��B!=/��İ"a�a�Ԡ�j��Ai�"f�7.YOy��y�� <�����׀�md�l(�'��BPcu�i�f��]��C%c��2���(��l�wx���N��U�|�Y������bK�
�Д�{��G���Ea�0�Q����I�Z�ތ�镸����� ���(��U�v�t�Y�Z�����-������#�M�oQ'gH�9ͳ c@�N���5M$���xE3qq#��t��x��&�I%���/�3��"UI�%E"�B\�f�A���Ec�Ӎ3��Z��$40��s*�j�N�����kN;'Ղ`�'h:cr���oo�H� ؅7y Ew>���}��aA�l-�)����>�J�r�����(W��a� 8*7tv}�t��v�f!_�y�TV��e�Al�揣�d~�Ri&���9S�s��j3�Y��8���(	���ga�`�.;�
����٦h�'�KA:F��Ύ�M��� ��M�y���Tn��C��q�W��B����)��)闾S�'�̇Ц%��X��4&|:Vfm��۝��ۀֹ�;X�4P]�א�c��D�Νy����P��bX�li�>���>RXcp�t��3_���,\#ӺꄥŻnj'd��`��"��c��� {����r��-�!��SE��#�5�A��{�u��;م8�Cl�ل��F*�y��	���"�I�p3�;�{��*]�.�*��W���_8� (���ƛu�H�s�*�S�'C��/%���z("�����'g�5�e��I�eG�#.,���WS�*ZC�\T֒�����W� ��� �ņ�D�|��H�9�Y��*S�`�*�������{��>(�֙@O4��*F����M��̵�t�U���JNB0"f@�" !�|{�f��K#�c��ߏx���C��s��ԡeLU����_
� `�p?q:�#I�V�>��Z2{�=-��u8@�J~j������p?���|	�A]V�ʲ5�V �ܴl�?Om�-�oV��%B�b_�����kE�7��t�>����4&��	��q�%al4-���6c2�m�n>��֊j��G�b��&�"b��~�� s�w #<|�P���&<#כW�`��У�7�����a�"+Ywj�g ZIGO|���7�nG�>�[�������ؚ�|���-yl{X8��/�c;�('\�1��ґ����*��[Z%h��d�)�ƀu�U�*Et��������c�R�v�?�F�0��[Ro株o�\G�2�@�u�:Yc����@��#�"���Q�ۀV68O��N//��p+�����Uj�-7�R�4 N�@�)�۔��ņݚ+>|l8�c���K�#x΍��/��V�����$��z��g-NF���!���ߊ�zY�����i
p�󃐾�V�#�������5,$��DX^�v߮wQ�\s��_��L�]cJ`Itf��DG����&[c[�� ���0�^*P��8|�Z�_l<�%��=�p�j\_�Ȣ�8�mJf����D!T����ͯl�q��G.$c�dS�������I�J�Qq^�P8�8V�@Ț�ײ��i8�� �<Lèh���?d�����޼�H1���$*��=�SrH��a��q���)Q�x8�`O*2�ڌ 6IR����U>�aX�����mgK��`�1><�n��$�+;Y=�at�lt�h�G]���gI���M�戱���l���)D���9�KAd�VƬ��=��)���ͧ}�x@�ܹ!Z��zc��ϐ	���-�7$v�/ye�n����^gX�����	�0޿�b�cX2!N�?�f�*G���C���4R�[r��i0DY
�C����-}̣��
��:˗������U��6+`V�B���ijg�Wh(E*Y��G}�#z.b�����5�7�ȭ&}��,Lx���ĢnD@�Jo��{N+׿���9�4�ah- +C�djp��)���%��i_+x�����?��x����.0�&]�/��K/��v��\I51a���AY��(4�j��ؖ }�#��)D��#�����w��ңT�H�>�^��#�����~T��ᅫlE�m� e�y}��3�����􄑨�hoe�s�?���9���*�q���&��Z�*�;^.���	��;��o��Ö8W �U#c)��G�̆$��-�,�����p����6��`UUxb��C��PI��mz(>HB��܊�}9�h�wģ�G8�lqfҙ�u�A�>�8�S��-���)5C�LA6�9Q��wD���O0i�����Gj�ut�)�����ʢ̓��n
���[�n�$��N�f�r- ����u����K|#�̡ ��=��Y�:<���Tf��qF!M�ajy�����y:~�-Ň?}�>��49��?^=�ö�8�z�tS��J����~C(�Y4��n��llP�8ٷ�g��ė>䉭[�%��F��7՗uTA/��ԧ�keDm�O!J����r��L��x���V���1��N��<w.�':A���aί�,I�^�6TC���ް��<^��/
4��o����y��0+d�7YZK���O5�����NԦ#o.cT�A�b{�Aw���k�%o�cKZ��\_�"j���@��r%J���]�ȷ��v��ƭ�i��˱'�+�Yq�0�FQ�8�2��1
�]�s�A1�����'��W�s��J��#���ΎF&3l��2"��>2:)q����>��!t۹�V�Mt�8��}>O�5����'H�Ch3��*��y�qW��rq�<���(A�Ǘ������Wz�� �l��5���M�����c�YbPH/'���������.�l��z�^�� ����'��\^���K6Y*�o<�w$�1 �(z�vX����Rz@|w�?/�2
�ll�a=5����Ho�c_�c��ZP5�d��>����Ɣ�73?g*rIܢX��u��-��z�����A��{J��ʺ�����txoڱaLw�/��������w��e�G(�1�[��W���jɬչN�!����M_j���lg�mHX�Ru7�H��e�l__X��K�aP�R�0F�����������)@s�U��J��hҞ��9�uF�ըI�,�B����l8M�8���k:ӑ�TD�N��CdOV� �>f�`I(�Y��n&sܟ8	�f2�GԷ�oTL4߉���|�s-�O��N���C� A�52T�	xА[9�T:Fѱ�ᱛ>�f	��D4ބ������-r��������:l,��kdk�>�[��ғ��8�"�\�s�<���1�Ԩ�6��6),����.�ՍWs���g�x�e�.����	/� ��$mg_�@wچ_&���w%!j�,��X��Lclۏg+��܂�h^����3h���{qy�͙��aR0��ج\��=-)^897D"�Bm 8Br�g����ޖ$��z��^�yj�1�[�H�rsa8�7#ļ��WU�\��@¶+��ط##�UQ�-X�R�>�����G8�r"q�|pZA~ǵ��9Zv�u�2��qdV�M>	�����5�F��HT4)~�ʮQr��
'�gj��nj��X*3��s�ժ��(e��jw�%�k��9dx�/�N'廓*WT��}�K!���$3�,P-n�bB�&�������i���%-a����6w�>��L��
b���UI�f�_���/tR'!b��O.ЗP��:ډ*O�d��EA�G6d��s$a��(䣪��Vor�	�F���'C�er�zb㯍�N�}1(<�[˱:�G�=:B��p.d�	3!������-v��g�VC$?]��Vyk�6Y1K�4�����{�QU�x���Rͤ��l
�SB
�y����ӵ=�9���N���z�HH/�\�l����,A���w�[�G��q�>{)j���P'@/��w�3}���\b�jH���Zi��%P�� z z�zZ$��(�� ;��� ������}z>��O�I�$�]q��f����L�Xf�Ӳ�#���>�	�Z�P+v69�����&|q�L��|E����n*=�L��]
�[c��
�PH����G�j�7�]�0�1~���Z���3߄ލ(}ͼl&������w/D�y��=z":�<�
��:\�S�\\>�@�f*�N��'ah�]��������sn�>����Ə'��!]�p�S��q��ʖ*�*w��뇱۞�!�>�Wk�k�;�A>Є�6X�7��Tд�Y�ܷ�O���$zT��9���������s�Y�`��xY�k���}��aՌ�P�"ؽ�|`$�F�����@��Q.*���H�E���<�&�$��ui�T��]-m�={�sY~��3ҧy��fINy~=w�Eᘛ�L,Z�?Ե�M��p�t�L�W];�dK4�>��ޅ���Y��X��m0�ٕаYܞp�6������_B��\�Іl��2�y�{m�f����^��t8�-�ϒ;ҏ�A��;�q�H�������@�)��m{�+����՚�2|M_�!�0&ɧ�E�aV�b����X��o"3,�sCD�>*�ۦ�L;�����SF+u}�9)}�o~�(�s@C�T�3[Ԭ����(s�n=JZ)m� �Oq�x;�/�{�Y#I&�<ڼ��&�ا�YӦ�b����3��#�0�!|���Hc/�������&y��04֏��db��v� O�5���+�{���o8�$qB�$N�u۵X�T�X
�r#��ȑ"�N">����v􋄏M�>�8�x'��%5�u�(bjS�bu ���`��?��q�ÿ ����V����\v�y��A� ��bl^��i�
�1�jS�U?�uoA���B��5�Q"�K/��HT�9������f�0���c�La8�gZx�p�{=�Rt���n��7�.�,�E�LU��	�o%�ܬ�[P!��&6_y��8��PIV��ϳh*��k}��n��@�na?��$���M"�0�N�X[�wn�z��Ȯ�A�" eQI�b]n)>�}��/�>2�A�I-f��:xzaB���$�A� ���4-�Z��e�8�ѡ��7��L6vh6��7��C,��;�"r�c��������0�m�\�mL�{ـ�X�?7qT/tN�U��<�� �Mg�c�?���d�pt}��xˢ��R
����g���U��	w�����?_�z$�R���� { �)+/6;������N� T�ji)����aq���@U��P5���viz��J+3�58�֣3.Q�#�_�x��j���:n��@[1���bS��^ϏPN�fBU��5k����2[�B5�LB�~
���`_ԏ3F�ӹ�ﺬn��U�)�(�;l�͆�n/N���&���Z�Y�����DN��]0:�����|�j"�]��V4�k��S_�����Mn�����I���K�>1�L����\�?�2��h�D�T���[J��7b�ƭM�~Q���#'~F`Ӝ/Z��5�I��i�� �)uB���p־i���ÉNZw��7�!��5F� ��1'�Y�d�ab(���V���!A��B�h��k\�cl�o���w��l�so�=�OFq�������6�DT!�X/W�Żo,;���F�
۬��֡<�vR^ZI淫wH	��[��q[�*?�Gt�{}�c�����SsIp����75A�ͺ�����v����_�W_rK��T	�͛���#�<p�c��Q���ǺUv�Y*f�y��X�\9uw�%/ٳ}3���^$ꏆ m��B��BO1*��8�Q@�5�q��[��)�w�~)�gD<����k��h�m��$k�^� ���|�����AO���8&�Z��{�@�9�I���$
���Z�dۊ�6ų[�T�J�y?F}|v�De��Ȋ�����0���q�ܩ�Yl�0Si:4��W�@�x5 ��#���ء�a�h��W=�%V��	�'�d7\��D�3��_2�9bˈ=rd���MA�4�
©�\���6��E�,bH8+���4��ӣ��w��>_0Q�!r��s�����x�D���b�����7ګU`���V�u��}
k��Kd�3<�E��,�����f�̅8+�����py��3��EU�]�Z�������=��;� �`f�Iu�WNŲy�����>�X��>��a ����fq|�-&0���~1dG����l�$�,�S �)b�𢁳�� �������E]�R4(�L �?�x7��	K�v�܎vs�` PD�����5���m"->-^�`�|K4��"��b��)):���gwmY�zF�Bڈr�!Ê�C�%!pnMŨ}�e�u�.cT�+\��e�Z���N2�"no���d�7�ی������
��N�ܤ�"`I�q�4qt�ғ	q�j�@m^��9{&?��A�ؒ(�����j�V�P(!5W��Az��b�����U"�/��F�� ��O�ŀ���\n/Ks�3����h싨�yh>�l9өK��{����̸�1K�uf���=�>xW�R�����k�	��sL'�[\]^����x8e�"��B����$u�����nc�@rr{��y�}�/���S�H��p͡�K���&T�.����}+����*@5�����#+��:�rأz{�5?iPEv���,\�̸�˄S���mL� �K������z��3��=eARd|��@%�#I.P����Q��j=����� �g��=���)*����g���l�2��=?Gd��4�:!��QK��o��*a�p��(p�xQ5b8�/��r0Ti��V��E��k����놸J�6�`,�p!e���睽3�mUĿ�\#�J���d|m�,�{$R��k��Dq{2��Jw	����Ə�Ͻ��@���?�GZ145�e�2��4N�M�����gs�;O�=�.Z�����e�ݫ���P*����32N����)��`+�g\����zis�����a�fz�$OC��6wMJ�ķ����|��av��@����^�e����(0A��"�����g�v�OX֤�%�՛��;L�?�$&QѤY�����_�a�)#��hғԨ<Pm˃f��KK�fk��xGh��0��!X-u��$>GDx5sg �V���^L��<�,^�%?C��.Q���n.]�	O���j��;]��1���)���{ u�u�?���k�;��WM�.,�����C���}��";]�y\�R>e&F2K�ߋ�Bq���zۡ4�K�/���P	����J�Ϧӵ�Q�"��kO�v��V�C��FH?k&o]{�A� ��ޭ�y��
c����4�޷4ꏭ�'.4ե��rU+���cz��W8ߗ����H2ϋ�E%��ѰY�~$$�Rc"�i���Z���t�(�cjU���-��8#�$������	�Y��W& F����l�����\�Wy�e��dמ��q�ѷ��3C����:6<���_�����Pĵ�\��}��F}8_~L��)��'|)�
�LVf�+��NRE�;a(K��.�+'�	��� PS��"=B���1�L�Ҟ�Ѣ�(��t���&��kf�iD���T��- -�9��'$Fn���0���Z����5�,u�ߊ1��P��%;��Yɴ���2��X��b$�$�ofW��C�i��מ�����r�R�]�)���ĻI/���e͊_�[��o�OD�PTh�:?O��jd5=��%� �0�5\�Z�g���^�1��̦^8���*E"�k}"��˞$��g� �]'OG|�d��ve�mB�X質�N�[���z���fn���8;z&��.s�؎��_��SE�f|�F������ƀP���>��.R���o�f2�^آ?�E�N��������LUr4�c��4�U��r��r�Y�kTV�R�]�mF��ѻ0�d����=�_iG0߼N[�º����>N�ݨ����ϼ��4t�o�-�M������~~����2I��D�ɉ��a0��p�b�*�،��12�BC\�y^�@$IW��sI�2�*�g��l�$\q'S�KA��8��t��;�V�$uݖ'%Yq���v�|��F1XK8&�̉��$IY��'�GI���'T�z�3u��z'*� F:�._K(��})�f�Q��)�L�k4�_�X%��Aı�&������I=�[���K6�%��B8�Ξ��>�N�س|)������`�}�� |�'N�`�L��}��K��ˢ��J� ����_$��8�*,���k9�:�^3�($�f�$�$Z�ƌ\�|��_�r�5Z������%^zNg���)�y��c>*���$gz�qv�C�ON8m̗����HJ�����3M��S�D�w�
u� �K�J��Th�$*rI>�RI�����v�AB�!�W�ŧ2+�,oj󾫼��5�}?�̂&�xA����F�o���G(�������H�t�+�T�4��P�$ӊ����n�Rh7�S���۸��q&Ƣcwl�a��-&aT�'t*Ǥ�EVZx��I���@�ɑ��� ^[#��%�ڒ|TJ�N1�P��2x�����>Oi86C��?�8f���/��.�:~@���Ԩ��|�&[�G3p=F�c�z� �S�S��/K���J���F2�����b�f%[�hvF�h�pdb:Z8���ܽ@2��c��7^��5�����U�{6�NsFH�LZ��g2w5�}e���/|5E����{D��9#s@F�4fԙ��Q~�K��<A��1���ܪ����d���_��,��6�U�\�j��?<�]+��K4�5����uA��Xx���;f(�b,m,pp��!I���ܩr�%�<��i�ܠ�����Y���"�G�M0���� �f�㱱c�������b���;;��fZ�ڠ��n!����R[Ya��{���1�L��Ha-�0Ĝ�#L�!��7�7H��d��w(��R}H�rm0ɑL���=^�I�3����1&�4�	�Z��ܮ���8����H/�:�i����5�5���a�/�\7z��.Ac��f�_ 0�c��@�&���3θiɗ��Q*-9>�l�"��J_�H��O���U�'p^qn��Ee�/�����Է{OD��mAori6LF���#V������ ��\d"%�"�=`��qҙ�	o�#ŷ��Y7(P�ܧ������Fӫ�����@b,P�kYq-�uP��dj��h���L)� ����DU���f�=X���q l�A�;) �L�����V��\rI�*�t�_"�6SH�C��E�h�p`�q�$��	j4 '���"��'x�B��v������|=��P�y���Ǜ����9vAz���H2�^xuh��XZi�6a�'��i� �b����^�f��~�:�����u���~Z@�#Y�͎��}��꘡�%io�N9��B�D%f�a�@:I��țw�I�3�eԶ4�3�%CA �b�ؠ�t��-Z�@�<����>s���(��v��,)}7@Y�4B�ľ0V�M�o#�d�2{0�#�	t�'�F ���+�<+�>*��Z=2�}fb�R���]0>;4����Oa��k4�7�
���9#��n��[x��ꢂ��H��q�Q^SWs1t�>��ԑ>�> �j��O��Xi���T�� �	%sǳDӅ?mC�Pޯ�;�a���Ha�Og�e8�Y�8��i$�~��l��|�Uf6��ͭV,װ�N������U�
-�S(�d(L����u\��-���6Ѳ�o8�����'��+����}&J���[��H��+�n��3��r�'2$�)k�i�K�lcF(����|�6����2��E�eh�e��<4u]���8QPun�oރ�F�$�YD�R����0e�t�I�ֹe���}ߝ�X��sXwN0ec
n�����
jqF$��	�k�� D�IP� N�ۓW�X���9U��R���*��Dvk��`�]��Ц?I{'X૵I��ۘ�������ʴ�zS��d]�9�Fֻ���@ ����ಕ�-"\z�G�Ds��P�y'&P[��bp�b�B�1�rT�d��g�׋��){�qdӣ�eM^����X1,MG>ݢ��5��4c=�]��z��ڈ�>6f�c���nP�z'�ȋ�w=5h����� ��5��C�>�(��!�i�7�����C$B��J�3x��n5�d	��ђ�a-���$�5�*{�Jf��w�ܵ�1ԽU�zd0欚)�%6M�T���cW� �~��o*طD`���;]�������5ljnJ�_�@����+/��;5<k��N����Q��"*��_�Zs�z]?K��s�p���K�S�!N٬`ȃ��%]�y�ì��+F�vԏ� X{��%'�<؅���f
���U&s;�c�{'�i����ф���g�K���,c�H3�\s3S��2�$:*���f��a%��=�|/��D�"��8��:��[7 \?j�G���a��F���i*��Mo#o��G� �bd� ���7�E����B(XߩR��q���
��~�D�)����d[���]wMKo)�Z�����tr�[0�G�\���'��,���d�NU�̞ \�X����Mu�<:9�4�C�����X���vn
�g�h�{�Ég�a�5/n�@���6���c���QW1]����p�sX���8�(k;(�"}w4�-T$�C�R�^k8�Y&i�5�EM����T$��;j?�����Vx�Q��6���,��&�� �9��ѯ��^#�����W.*s���~�jQ��f)P�la;�!ѩ�����f08����$3������7������������u���3���lUC����C���@�>���H栗.D���kXNY�����ƚVo`�@^At��w�Ͻ�u���8��˲�)�5����k����7�� x�{�+�	$��j�E��ҪE��kG-����`�(BQ�'���B�̬5�Wr9EM�ښ�oR���`Zj��qeA�ÉI|,�ڴi��j��ѐ���4Qgn�D���ݧn4�!߼^�rA�"�,f����ok��'��nE3�*.�=���#�2Yw�y������Ng�;��f�@���LU)�D�[�(�oxD(�'�|]�^�&۬���\���-Qr�^�9@��ؑ|�Ϩ*��|�}�kr=����M��&Ѐ��@VA���� �Զ�r�aY��C���$'��RKZ����4�_@E)�rH�/�L6�]���u�8 �[�.(  ��߄Y�iz��	�l�4y��i�*zi�d"��spA@{3���e�T��v�d�^���@�\D��>L�� ��Ѡ����.ү63���r'aϽ{k��h�ȱ�^��W�lh�ߥ������'"q�Ŏr#�CdU�V6�(+��DB�����?�\X�غp�50�6�J�Y6U���͛�=����W��E�%R��*ՏZG��FP#b�Gs�I/��X_��c�U˔�� �5��4��[���=q&��)�ɞmc�gؠH��y7��߈ʋ�e ����ֽm�]J�%o1�w�@-wN;��3-���e�z���� }3�v9����5��3|�7����3J��}2Y���zb%ļ�;`�����zR
�������m��;Һ���󍼓��+���@���Q���N\��9-
�7�Qƒ������E"��l���E%R8lݍ�\�큖ӑF`c�{�������K���߇��,�����x�v���iܯ���ky+�`0��c?���ڇWq�p��iD�0��=p��s���F���A��Ϳ���#s�p�.�heAQ���[Ģ��{/���� �?��Ƽ�݆B&�lJ�ev�/�P@)�c)�]�����w2��ı�\�-�)V�r�OlxBu���3����׃v����u��*Y�V�"����s�I��N����h����]{��p� �Q+/�)��9�s��_�.�Ë7ԌUV7G�) �m󙲚q�b����2�[WX�f�:/�G�Z�_���Ƀ�v\Rz�Vl���k����>a[��3�$N�X��L䞃��4���9r��Y[oZڛ�{��eG	�{r�!ز� ��&���۞`�ܗf"��!4>i�9��.��"�9��S�D���l����S���(�(vMF]%sۙ�,W�O��#@�:����`��5��(m�=@��&��b547y��:�kBˊ��ۨk�sy��݋� ��T���ۧXs��(��T�ߋ�����"�)�y#��k��BY:g�����Sd������2�	N�7in�wld.�@�pp�'ҐN��5D��ۅD�s=)���[�h* `�'�.���sԸ�L]Dy��e<�A@ӫvƷ��r��2�M�{���g�|�z�n[��],`�����6�?	�ҫ�;*WK�Ɓ��M/_���^������c�-���ϯ�r5&Z
��x���^�b]A�������[�Ho*�����E����{���c�h��ӹ�Q���ޑ��b_b�r���Fh-^;sD������1�����­�C��zjg�gyΐ���b�8�%�tv��s���s���YX�1�^w=3�4�����*xĪ�%6L������d(tYl�2�c�k���}�sg�-'��s�*$�����G
?�,Tx�d�^,Gp��p�i��$�ix��絯u���o%�NRi/��c���noڷ�/��t]hI��c\�<���*�z��/��!�P6�k�"�byJ���cL��#5Rh&f��n�y��*�%{�l�����P���rx=a���~�	s�eH���Y���`�?�yC���[���X��o�U�Y&!N�*�4������-[ج��S(z6��|�Fa���ql��
��M�.�#�
\�_�n�U@�EX߰[��ߧʨ逍(6�,S� o�<���'�F N(,y��-ҽ_\�L.���h�)eΈ��o�\I��M��.:X:b�V=��?krjgU����l鹔R*I�H\R�kãܣ󥖮v3��K��C�ԁ!2��F�s'��C��m��3xdI��%�MB\�g��imr{��a`8vahM6��%����g��<dƇ�ٝR�C��V�{�G�
�%���TN�p�B�c���Rӈh��򴚱�h]`�^^�c�v����>��/�"��ǀ;��� �!�c#rtL��Gdd�6Ck4�5���$9�;d�漀�|y-��3��J�YPs����[�eJ�'�)��k�p�>H6キe�˘,T�����,E!_;*�0��H�ZZ���Gi�$✣�kt�?��WD�I»�L�[助_�?E�_4�dp��u1�ƈI����m�Z$�$`�[����P��xTC?�'���>T�t8[>cM.ܗ�
��g?A�W��#.�2��o$��}a��+(��1��wϣ5x�˩��z�&���vlsЁ>$�&(ݖl!��T��� 4�@RRGEϘd�O@��<�p�	�%�L�7O�\��U4Hp�[�����H>ug=,�2>�T���@l�$�c�W�Z�v�Zd���F�uB������?9���h 5�W㋯�^��5����GNh����,�����ċZ5z��>EXJ�p��d�e�����?�jy�����¯���n*|��+!�n�q�*,��O�J��v{%�m�\�����=Ho��fN^hh}���3�r�g�a���G'K/�8�%p
�u�r���0��2(-���4�p%��O2��;�q��ڋ�^��l[+�%�/�I���9�0�gu�ln�v\��g4�dћiϽfb�K���B3����:�>J�"y��[vሃ�Hʒܙg����I�/>��L^v���ߛ�|6屠>�\����i�y�E(,60v3qLAb��i��,�΂�1<>�1�`I�&�eǔ�z{+�R�rUFܩ�&E�>���:.i���&�y�k/���\�/݈ .��u��1��3���LBW��+�;�@(�n��m����oO~��yҜ���f���&�Oʞ0�������L؜F6�$���V�Pq0y���o�a|���K{��2�?o�d7�����&��Od��ք7`w?��T<+�:�\"hG@�(m�rj������e~[���@x�f;!��d��w�G2���W��jlr����Ͽ_=v�)j��p���?H�m�u1#��d�g��Kfra��xˬ@���/넌�U�d���v�����{���G�p&+�����)���\G�1�` *]U�/�u���V�$o���5��S�$&좺�^.�"�wO�N�j���L�U+&UC�e�Х(c���V4����n�X����7�x�K�a�_g�p+q���g�y���s�z�L��V�	O�U���6�F�S]���ZBVc��Q ٞ
���g�WWJyd�����	xb>`�"8	;�����2
�\�����.;,�P!�3���G�+!������r�N����R����!bf���d2�0KG%�N7�Dm��.�0��l�r<_~���5��ŷ
/c��6��Z(���/7~'>���]������Ϻ���rB.���*c������?]�����Z�&#M�[]���� 7IL��ʷs���5a�=�4P#������br,b?	m'�q+�K��
�S��	�{�*��	�-�XKx����6 [h _���H������� ���ol���!`I�7�|@WW�crȐ s�@J�Ø�L4�Q����#��k�D�M흔bs4A���LU ?�+�n�����W��Q��ްH�M,�0���;%j�d�T��n����׼��ά�S	7Q�c1d�X��mS?�muW*M�20�W;/�!aW�|07�	sͨ�f��/��A��W���/�)��j��}Y�s���c.�J��S�>����&�����ޅJ��G��1N H��[t�wU!+{���Y�?��a�΁,Z�]|=*n��ؚs^�b�>Ƕ��_����s HM�����WIV�e6	��[��ʧ��͌;�k֙�1��6�/<�p����,�ڲ�1���Y�R~Cx���jR��ݸ���?=2<m@n�����X�R�w����R>���z�[#*��K�)��x
t���-@m_;-���b�\�c;���í���q�nJ85#�i��������m�yæܽ���P����bڍT���k�7Q�;�8Pn:I������pwJ?>�S�OU͌�ZF���iH���ېѯ���B���߇����ɔ �(ܝ6*5��x�V}�.�9������3������j.Y���#���0�ǵ��*:�|���$u�ݭ+���O�+O��������G�?�~���p�f�DE����Z���"W����j�u�9��M �3�0��z�,1-��&B �r�ݮđC�T�"��?�qZI�8���V�>"��.i��N�=HE��� ��e��H�,�|�AE�o8��c�LWoZl?��6���j�Y��uH[��	�۩a���-�FI���F��3�z��
�1�i�4BD&�mca�0vme8��5����B�m��.���LQ�(�W8���@O;��p�Nl�{,`��U�vT�֚�p����u�L�R#Ia���5'�@�snC��JIz����?��P퐥O2q ����"�vD�7W�� �|k��d����pf�mj}3i��UQ�σ~���dgm���)^�k�g�H2m�B����Dj�_}�Ci��MN;�$R�ȲG~�Ƭ3p����][��-l�	�(� �Lޘ���!�D�+dL��5�E ����Dٝ�,eĺ+���ċ�y�F���yY�Eų������R�opG�$���wu�����팪�mV�����RE�����s��6Cȁ>d��r� }ާ��I��a�@�;9K%��@̄~�o�
̤t��P��Y�: �k����n�{�sj��(���z���o,�_�	�����O�#����m7�a�%��2���C��A~�B�|������ӹ�ǵyO�LCf��aq��|�#ޖi!�{"!�<}Z�?#A�/������R�rRR���2����],��5�-�7�J���V��.V��(4�cy�C|��K{����_�7��?̭7���0J��M�j �T�|�I~�<֛��}|~a��ճ�W�B��?[�EUF���f�����1l�Bh���9��z��]�GF
��vV�c�*�q����m��5�H�x����Z��WQ�!��840�yeG��w���"���ӭ5R�ъߺ7ad�U{c �����=f����w+pD� ,�5΋�i�w�C�`Pn��;�e�7�_��5]��V>�f�D�e^DD� ����͔^�ڔ_���
��Pw�.�hV�����g>�ʱ�"|�Rq�ʸ�uN���%��q��ȱ��scM'cS
��N]��M�3{���t"D|�E�m�=���B���G�\K�p��an���fȯ`]�V�%Z呾�+1j/(YV�uR���mQa�N�CGg��Pm�L�)]��J�}V��._�_d��Xב��G!%s���i���VBkkV) T�o�ڥ��ť�h͈��@�J7P��s���=�/$���*�B@��;,v_<X�L�z���+Z�ڋ�*�,2�WCf~�7�5c�K��UU�I>f�f���W����v�/X x ��eM&H��dQ˫W��!��Z��ʾ�m7e+���d��zGypյ�E�3��z�k
�^��Ok�GR�9k�)L��dp.Z#�;f�RU���*�{���~!���z������<Q!�ϛ�#[�w�Ә�>uL�U��Q�.T�1(9J˼�_��3���1�$�T��8b�ܻ�6��-*{��(��	Q����҉̒z��q�0�8�8�b�+�-[�� ��&�������]��^l�T��[�V��Ӡ��R���7P�-�.!l{d<�M�:��׳U�I��Wd�M�<g�]�$�Ƙ�����C��0��{V V�kZ��2hfU��A+uR�n[�A��D�����m9��em<����|`>�u^��m��X���ܛ��O�\�K�e�lĶ��ԙ�@g ��ku5 �D�0��������=�����qۥF���(����<6�a�ߌ�
������*Ӗ����:]joB�6�BH�cR�	8Z|�Ú�D!q�u^B�;��!�$��PY�����~�~�ڳ1=����	��Ż�������L�̮��H̱���}��o��I/��J{1��C=�*���qf�E�C�^��a��?���Ff�Li��U�*l~�=jJ6��-4T�K��d��(�	�y�J+�f�N��i,�S�He5��7\����\�[X[�*6�3��ߕq	�~����@���'�ŉQ��� cZGM�L��5g�H~�q���@��:JBH��)���-��Ud���ɡ���>��Y,�'��	�'u#֦-v��T23L9�)!�$+elvN:cE�$b:\v��P���W�����@�}������(����lr�?C��g!�����5�Ñ@"��O�Z��G�P:�C�+��+�]"� ����кq��2�K��_{����9��`/�(�����da�㰃$��� ^�)F݆�p�`Q�t���)�g�CS$��*�}9IF�Xe�gO�TO7�iޚv&�+�4M�ok�q�6��Do�( qP��%E�2|�jV|1 �^�Z%���(u��N6��'9p���=��S�N�ƹ10��l?4Ka�*m�X���.N��{�v�s��]Հ�z`��q������jl�0���D�b���5���>�XxDp���z�3s�b?�e��<�-T�sZ�|������+1@XLh�:���R�ܽ��6��G��[#�v�u��4	�R��/�����W�ݹ>�-Xָ_ú����v#�]}s:� z7r
�e�~Vn��>V:��8�R���Ւ�	��_�.��&;r��l5�3�w����	.�N6�;�������"4F<݌�	�� �?�K(�>�T`K�30V��;�n�����"�<)�q?�U
�D{���dv׵�#�}����;:S�DXme�h_i�19_ (�W��ic�@�*�=w��~��������cya����>�z�4�`YX3e����B�Y�n��xf��U�P��,�݀�K5��k8�2PY�:�t��	����{���Z1y�������3m35�n��c��J�i���I�z�R7gz����"��8�w�V<W��,G�(�r������Y��� ~�A��w�Ճ�W���l,'�n�}�������nw��O����Ҡۓb�E����s��j��T�^��n��lزF$�R�B��e#��u�Ƙ�Ԁ�V���if����8<�`ҭ���w\G �?��+|�=.�q��-�D�8��]���eN�/{����A����uJG=���Jb%\�q
|\�sʩGds:�t�na 7�4�Z�]�A�##0f�  ���	k��޶�J��1ln��Ȼ�Y/��k�̴����5�'ܸ �%b)�G�o.� �&���hd�Q���94]k�I,�Ɉ��PbV͜pJ��\#����0H�,D��YP��W=<HX@/n(O��X��l�sPYE�!����ؖ��[M��b'Q������T�~��
�U>�6"l�7��ZŃ��H)��QE��4�0�&�.�	�@4ڈ�	Wl�:R(�^¤ћo[�	���=B���Z��q�h0�?�2�?6��Qqr�7�'���E��&2B���r��0�������>x��GĬ�Ri�OSz��=a�����>�����a�r/���鲪��e�,2Aãn�H��������I)p��k�S�KA�_�������B�;l�v�{�q!����c�Ux۴�D.e�>$�|�[wi���5To����2#!遜0,�� /x��$��=f�Zt��@�6. 5V�Ո]�0�Y�N�����j>w�q��Ӄp)���>���+�Ȏg�8��"�bPٚC��3���4ѐ�����k~O�$f�<Si�]8��X��F������*�v(�nzhO�0��f��9����ߏ����#�&�W��'5�ٗ<a���l{s�5�C��tO��&�ܴ=?P=�A�a��l"��ɣ
q���q��R1��nP?P6H �)�4���Qp&cH���o��������n�X�DC�$o�%,O��*xMڼ��ψ��W�����!N%�[���,���*�d�f�E�(���Jk餞 ~�xb��\t��ƭVʃ�b.���s��_�amC<[V�P<넡<��kk?��^;y|��~��j�:(u�����z?-5���9�(�A�o��/����e�k�{�~����y��ٴ�1Sޑ;��h���������`5Ӈp~4���R
k��YG]�E�*�n�&�D�UĂ�VQ��r�J��q��O����+h�v	L��y��>A;%�a�Bך��>g� DWٛW��py.f��F+}����j�ۀ�Վn�������9�h����� ����Ė]�gE��9_D��H��j3�q�2�V1����6>%QS�)?�;��~+��;��Ӈ[�RQ2�׆ҌE����
`0ӓ�s9�#	�i�`�kj�>$� Ćzf��l��1��J�FL-�]����d:��KEtWsm��N��aXNU���2Gچ�c���&��K��7��AI�c�4 G���V����L�+��c&@��W�_�o�F�����)'m�F�`3��C�U�h�DE��e?g\Js#�u�\�^���/�փ��������f�y�+P�2{�K'z�*n���2���������V&4����f��������
�e��Od4/@{��T	���gE�#������o�G�*��v���(�o;��j]�^�x#��eL�w��]0�==u-!���/	��?BM��cH��30�X�����/�c鯷� �Pq���/]dHr	ϴ�1>�Z-���h���	C��ҷ�+�e.غ�M�d�Fmi:��թ�h���U\qE[�~FA{����\��M�{-�c�a:ƻaS��;�������EX#i����Nm��ΐ� 6�d�h>�S���}�>��>�T�����oB�Ƕ���\bmu�i�]�.�by�V=Ґ��W}��0�I:[4��_(_ؕǇj_� �l��SBQ�#	��[Yb�` x:�/a{��/:���R^>�My��Sʻ��S�
S�?����y�����?t�]��x �:���Z�i.�f�"1jF:|��0B<F����OS������L�;��IH��)KԬ��Qn$��)b�Vz�� A�Q9���eX|B�n�/��F�������˰A��B��-�pi����ä�st�ٴ.������U�} �dQz�-�u���d�y�_Mx� gRƪ����+���
o�e~�n��l͍���[��o�J�p�FqǱZ#9�Pt�&|��<$\g���� D%J%���e �+; �r���TѮ�e�ɗػ9}�q�����=g�F�}�O���h��"�>���B�����3C0���~e��z[>�&������H&12ب_�P���5R˞��9{^d�}����&�z���RH��`���q��^�/�ur��S����P��c��2��l�nWd-�L�bg},O��8��5�.����]��_{�f"���F
j+��V����;�yA�/��d�U������z���t��(ff�:U�2�s���:M���0�u8.���{Y	s�"|���:x����ӓs}�ȵǵ��JCH@���_��7y��;W7R6Z�
��)C�:�^�LsJ�ۈt,ˊ�ugT���olWm��sN@�P�2	V���\��ә��w����?��( fi�ʪ�Bq�[3���}Ѐrc&�c"���y�py?�j޿��zߒ5�� S��H[iXw��\j�mO��M�Z��&s�D�T���n���K}���:5�b��M�G��a���L'���8��
c�l����5�*E@Y�:s���XQ� K����� �'�+��7�J���#��Aj9��D�F����h�}]�tP�D_�9��'骣��3���}��,�֎�> ��8��A+���$G��]3���W��j��G:��)w�� �θ��{�0Q+��<�ؽs�k=6!�E��v-�6ߦ�ϼ�I�+�_,�i���ׇ�*6����y�͡�p;���7""e�9`d�)RA����w���ޑ�$��:���}ӂ#����u���<��|]M��U��4zUY����[
���q�{9�r@>��M'X���w�3nMԜ979
�H3��`!�l/�C n��}~M֒<���8'O�J[�&��R�+��?{i�$�E11�٬߲���vO�Ϙy��[kH�Mo�h�?A�HA���K>�~
�O�FD$���f�R(���W��7�i6�Js��3�ߎ<���T�Ď�"�}�[���	_����札m��/��rSp�0?��U6$�Q�!�����6J���^���!�ù�����,(,�8�YԤ��&�ދ��Z����-|U���H[�H��g���]ŏ�q!M� C�4��ӓ�=�J�`6w�ݴ|��r���'W��>\���I�t䄁��k+�e�~�.ONU�~�Ԕ�<'�>H���p��?�j+fI]�0=�P9#�0�Gߕ$��SL<d��?�ё�
 !t�}}��Hy#�">ݭ���&�T8�*�߈�����!/��QrKZ���&y�|>�.!x���CE�.��^#��Z��#7�>�7��IA.��:
��Q�y�A�X�6Y�v�&�D����~��p�K	D�N9G&����톰�G��d�͡�g�k?)�Y*x����@�?v*hZ]����2���'s���`Y\)>)I���7�y�����I�{y��y���'��!�ҙ�4*~ l1H���~��ڝhg��}����$���
�D�P�ܧZ�'��6�Aڿ����Hm\Y��"�[#D���0�� �ãֈ�b�薉Á�M��n5�2���塿���t��.#����*t]�L8�rn*��T��x�҉ñ�.�~�I}0�h��3=��jl9�Qp��&��`��]�$���xc5�z����@���)�~(�Qu��BĢZ`}b�7[/��k�� VK��@��#����z{C��(����E���Ð����LW��~�JtVvA�$	��A*y��qb)A��VT3"o	Eَ�)H/lBs�bܙ+:��Djs|� Jdi��}��+U������9�Cj�K�_�:*��LW��>۟�w:�2O�����<IgӓTt�"���0h|��q���K84 ����wj��`��s?�
��
Ҕs �F:M��.8����+�үfxzg�8PAl���P`�9������s��?m#qړ�FH��������"�[c�m"�6���E�!��~��Lz�rg�N�]j�db�U�a��A!K(.YtU������`|�Avz�:h�rs�F7e��J��Y�ܦ����NR 1
�_��4��2�}Z���d.�K#�3<y�m�� �H��F/���U�~�{�T?�S�\�:Fxg2WL����L�>�'\[W4<� �5��.��(z0Xe,��vE��u��$D�o~�H-׻#��)<�HǞx2-���Lq2��Y��{���z!�}Ն�����<@� �]���&�}���rW�ŦQ53<�_�������F|H�f���~��1�zN��k_�ګܚ��R�����Ѩ�Vhc������������=��2���ʺ����~m�L��E��)������7�>���W&d��b���c-�|��H�O�ӥA�����Z������x!0�7�����>uD�y�����xm�����} 8��)��)2}JƬ�QV��[��l��s����vH!�
h�U\X1�6ӂ��_��qCb=ώ��1#h+�;��$�}3�;^� H�[0Gx�X�PA���.[ى�Mmǒ���� g1^w��h�5�c���w���
��� V���]HܶZ㕾���������Hbd��"U.W�*Ϣ�8�5;l�L�a���-ӏ�O�R��8e�@r�+�Pȼ�@��tݧ�Nv�pv���k� �f���+�}��AV��z�1O��ο��º�u��!P!*0�@�ል�h��o�؂qA/&��o	^jM`�a�;���F���rX�od2�Pz��̢�&��-2��F5�[�6�Ȝ�5_��;�.��WX�9�4�/D�![�0z�J1�OH)��\C�ܲ�N��m�k)Ёr����H���z"��:-��l|�����c׻0��'��,��@=+���C|��X���i*�Ny�֤�h������Z8�qu�� ŲMj͝��'A
L�MA�y2����n
�s��1�Q�JE��b���e�&�f�U$�Y�Z�q9��0�<�Ѣ�� �/���	�z�77 �����p���ͺi^���:8�HVpr[��Ԙ��hR�v��"��� ^�d'�0t�B$fz�!d���p�o�ޢ3�^�ڵ�D4w�4���VxP�$�9�Y���Zt$���|ܗ����D^#s��;��ڱ�1E�-@���8�F
�g��D�}~��ɐ*1a�1q<�pV��Je����J��[��=��ݵA^�]�^Ӿn4�AjB�'�!/�b�2]�C; ҾV���M��n��cv����İ�]�fذ��G�#�;D'�Y"��;�Me�Wby��b� ��x�Z ��ޣ��4�i�?&4�	(3�h���
�
B���袜��ZaEw:�����¹ƔE�@���0���Fd>��$�\��Fyx*ޟ ��u�]�<<P� q�O�X��@���>�KF �сCTZ7�U'_��EnC�ݤ��T�8��4�;;h
�ƈ�ҳ�i�?��sHڙV�y�8TSy���
�	+��v����ysOx�B��[�+[Z2�����n�s�8��M+���瑙jƓ1h�O
R�����Jr�b����.3��>��M�6��CE��,�qy짱-!����+���Y�]��Ě��U](�b�&���X�A����Կt�U	�O��i�}E��2�I(L�G�b�����ѡ|�O�G���Q6л�׆;��/׉{�!�t�!�n�x3	\+�G`𮲉�M���QWOO����hJ����k%`�]<�9��J�� �r�-���fL<�J]>�:��\��*�Ĉtg��h�7`�!z�� \�l�x��uS���^2�$����&�u��	�_�BD8�n�LAW�7ű����l����ރ���\K��M����
:%����oX��rUf�{�tz�c�v���cw�/a�3����[�n�����\�������J��jԢ�j4�10\s�YFjD��r���;�Y��ˑҷ�Y����nj�������s:� �9W��A������wJ���3�?���`�k�r�ډ	�Xa��Рx��ޢs���glT�bQ�N�Y9��;x���?V�� �����0h2��V;1mA��ͦ�,����E(ۛ�U��#��.r�Pvذ3�3b�3˧�����H��Toh�LJ����_�S��K@�����'pF�kq���G�����=�\ɩ���f^6���pt��Ժ�����1�����t�"��Q70{z�s2��%����d�Y�LE���p���r�Ns�R������*[� ��7��N����������B$����ǺhUIqz�Z[�D�>�-�oO�l�ɋv�f4��S�(�������)
�#���L��^k�B�_^D�C˜�������_[���=��~b�-.��X߳/��c�3 ����`qH�өU��T�| )�9�-C����V��{��Ħ�(H����פ��[q��{M��\ H�B?��2��Q6�X8�Nf�d���<�|��c��H�\3���F4;K���ȐD��8���TD��5^x�4=Zf��'�ʉn���X!��0EP�ʧ�h�θ�����q%Ɖ@�jT�tCX�<���T�=�q38���G�j�SQlcU�v�zG؆�5 ����Y��F��B��T]���j�:a�&EL���n'r��D�J\�Y,���9��d���$drz�wY���t��5��l��sJ���+����\е:���Q��H���_fĭ|�5dM`X��Yr�E$��U�M�e�ړeÃ|��C ��$&�'�W䀛����u�?��&:�6�i���9�jeӭ��/��Er�ί�+�lrX�Dn�t�ͩ���?!'���vb���� �U�A�E-�Odx�O%Joyj��X�`���oX'�r�q�^<�m�Xg{?y�m�	B����&r&ouN/�DU���D��T���\���I�8�|!�l�����%tֵu9S��jrBYL�I � �y��݂��uTf�?)�Om����6�-=��Bg9A_5�� �JkO�	E�u2�����L$���C��� fy��h�����u1 kNy�,#��#\�$`6.�k�k��4�\��޲Ƃ|��D�N���,$KA>˟�nKO���f���nꇟ��0�H��7�
n�����?�v���AV�YI]�w�H���ς��n��^)x��t4��5^���rT�F�=U����m���C��'�~z�#��K��jd@���}�)�ա�`�x�U9�(T��$~G�r<�>���!K�C}�I��ϝA >�s^R;�珩R6S���L�3�T����3uם��^ɀqGo�E=6���H�9� �������ș]D1�!��7�>g��!�}K/�<E�Gq9�o"q�p��p�$�>K�
���{������[)RV�L�;B�6�[*����س���i���̝}�g�DZ���G�=)������'�sm�kx���j�f�x`_���2�oqV�-�sI1a�v"Z(�=�[
���[tV�Cv����ġ�ƒl�~�/=ƻ��5�n�AQ~�W2��r����:'&�rv�Ͽw��h-m#��#Ls�����`"� �M�6O��9��`hOA]��i����l�XA�BtnW���?K+/ ��j=I�ƶe���s��-��/�k<����<��G���	�civ� Z��@Nk)��<��E�QȏT+fc��'��	�5'XL��j���<ف���%36�l�����n��J2��0PH�p����"E�� ��q�{�8�-���0���E����j����CH�J)3��N4�SO�a������K�)�i�9���:m4+ m���o1%�7{լ����C��fڮ�3���[����~)��N�Ha#bR�*��$CX�L�C�k�0�~+-�^�/}�k]�Yv�BX���{?bp%�c$��ѿ�F���*��i�E�3��d��\/A�8�+S��ّ����A�w�T�TcZ�g�&_l{�Z)ַ��Jn�͠?�)�]���]ɲE|J��=]����6E�&ZE4�&i2;P��7߲L��#<8O+&�
|��O�^��B��������Ϟ�&uFj��:�,5QU��0�RL�y���I,S�pS^��u��M+�h�Ya;`9�g8�����IV:��u2���tKc^{������W:Cwa�O����+6���Q�`���QlA9,�v�5T�3�L��ּjL4^q��u��~2ҲImT�*�N؜>�ҐY�Ht���g��T|��rw@��%�dV��7�N��\�\,Ԝu>u6l3w��fX��qS��+N'���<���aM&lQ`=�a��#K&W�'�I�S�gI�bP�J[���#p�i�o\�N���N�N����
�� �cw �Y0`Ťș���� ��_p��줋��k�B3ت�q��r�\ILL���U��#7�_�?70٭��3��wI�R���+�9�Dm�������}Kb��� e��%�w`aնL(8��k�70ݖ�D�(1 �S9F��R�5X���x��n++;��X)�bET0L����J2o�fOr{��`�=����Z���g�vt�"}�g�h�Z����e^^�N@����RQ���UH���(Gݍ�!�?Hmm�0�``�tY�n{T	�P�I�c�<:�t ������qU�܊�lA�l�-%v�����9�D�=��	���Z[���F���Ϭ�MW�K���(�jwv-!{h��
g�\����g�*��Ӟ��<B�)W��y�*@Z�39�8����+�^	�\횠��8�B`0��\6�����L25��r�k�k|u+�E�U�A�_���|9�Ѽ	��Rd�!�Kp1�,j�Ó��EF�2�K���1Q�<����,A���sku#V?���6����_���$d���"(��n$a�qE�vy�Y)w�Y�M0�(��]��JQ�y��-��V8s�©�=#�9���>�l�/���Kz�+:���HO1�R��V�
0l���L��""�#�-�8��cEU�\b����]��y�	&~�B����E�*�͊�f���.\&��6��t�n%<u?�"3-���W�,H]�$��}��+��M������p�%}WtN��N�T<>Z��X
�����{G�7�q�'93p��\����F<DJ�	,ߤ��'x�A <���̰���@�c�X�s�q�h
��j�T]vrߪ��ގ
��ЙD#5o���^e������k�¶�m�u��|���XI؋�k��X��9�|}���<���*R��g�aP�V�l���s�2363uFZ�M�ٶ�ˮA��� !E���D.�~te�n?��	�Ե�z{%�y#������#�t�Y�p.�ڳ�j~Y6����/�z�4�T|�Kw�A���7��M����C��So��D�1|�8PP�KtbXy�	{����3� �������暥1�8<��8%k�?Y"�&3�#���󭄸T��B�LA,�3���w�g(q�f0�/:1�" PaqYkd*-С3�q3�q��'������f ��^�h�m81���5F~�O��rM
;�8��Ĉ�Di�3P�ɉ2�P�"�C�^=��"\���D~�C��ɇ�3����q��
fd]��7� P���w������Ջ4L�%��!@a�$xʷ[�E`ph�X*�|���k_	Xc�O�:Ŏ�Up��Zi��Y�6b�qe���m�2�\/�r�_Es����dX�`��	�+�j��`]@����Z�J���zB��m�]I�$�z97JP��?�ptW,F��3�h�;����94���&Ai*iz�g��K��)����Q����4�$%������-���h��e��j�ܺ���&�h����2�)��7�N%�cd~D�-DR�[��{ko�
mc{�P-��B!��Wx|@�[�iW�߀]�T�C���J��i�k�鹽�dO��TcDy��i�ЈE���CD�=��@�u(Bq���{�:D�u���K�*3�߾2��ue;��P����A�p�p_�A�v��P��g�Ӳ9*[|�X�����^�˙��r�r>��hre��{��p�84��GL�b���]/S$$�=���r	7J���&_��uO� 7x����s�M��`1F~�S9[����2����}�ӏX @_p-fw���7�ϗf�X��d���G��at�t�R��ɫ�ڨ6�v�C$ �s|�H���0�"��!���=f�F�%�)�b����Wc��(!�cw����U�� ��QJ��{)�.�(���:܎�4�eU�ST��O��2���h�P����h�qԸ!O�N= �@�����NP�-���}h��㻒�r�j�o�p:2���^
�s�jJ�Z�̯�R��E��1'�?ⲯ�h-��3'�[1(�/j�M�KPO�P6�c�f�pz	�f�u(����O<ʓ�ʙ�2���vC�̂��s>���[:�\�j�	2w���|L�.t��h;Xg��T(C���
���+K�!�af��$��ad~��[���vU9<�Rrc�>�>Ș���P���)k٫dg�Rc���gK��Ud��LR�����J�p��װr���JNԍop�����P��H�@"���	�hm��|܂'Hh��o��VM�}���<i�=V�&����t��Q���:��,�v��M���A@�s�Rs9^RYݳ��@Ry����i��̸��]�jk��߷��"�S��e��h]9���&Mºd���w/�ŅoY���%����%�X�����;lJ����J�jY���-T0iOvq�g����x��}�k������G�`���-O�B'�T�8=���!�I&�ID�X{F��f�4|Aq�o#��o�:�f��7�R������\A�np�k)�
JX&7�V�ºNf)���ʹ!����-�U-F7`�(�&�E%����耪���LL�o�K�A�w��4�\n�[^_֩���K����;&���Y�ƯW�����F~��-l����b��#�>��]E�z�u�4�v�L�;�-�c�Q�7c/Վ�I4-5�_-PƍSMN�J[��t�Zc{����މY�:��g_��8��u��~Y��{�	2��(�� ��HȝU�'<����l�ї�NgX� � ��7�V�G'w��D�����:3/Y��Y�_d����"�5��;u��,dOৗxRxx���Q�R?I��mq �|5�YxC��:j	��<^�"��Kݜ�L�2 0�ّ�4���e�7=������3�_�m@�{�Q���ANc�Sᶦ��M���R���Ps���1v��!���v��>��f��.T� Y�r����xa��H�z{��b^���ۼNI*�'>Q
ń��LqiΈ�h��\_��APy��qWj��g�n�Lv��f�ܤ�Q台��}���W��B���$}Ck0L�U��B�¯�;��#A�nMH	 �,��8Szkl�2��:~" %B���)u:үtz!ln)#r,]�B;T�� ��L7F�
�#~@G��
�J�X5o�f@��0���Vw�� �3��ui�̘v�A�����6�����a��M?}en!&BաX�m�_���$��\�;D-�<TQ^����N��J ���j%�#�iuƺ���Z�t&���}6�d��$�L�w���rD����Q�i�ר8h433qqV�B�@ē2���b�XG�]�Ibp��_l��F���М��]��j��X4�'��!Xb�$\��!��{�_�cя�A���$UC�1�w�]b���؎:v�^+��4�=G�4i�c�܏����i�a�AZ~����q���}	SG�{�f���>
��l��Lr�\�3��{�|@�\b�RR|�ͽ ��-�*��#~�0������ɵ�A>��C����?�3��tg%��V���w��4��~f}�R'Ȓŋ)����:~r�{�hI�b��&����:�Y���F��`�%Z�O��<��7[������yl�C��z�xFř���� gn	�	�B9R-˕��r��tKc�̵ky�E�wmz-C]�ב\v�B1~Du=
9�s���q�ÒR�BPo���]<69�9���E�K��D��˴��8'�qpE�����1����T �kX�׃\���E~{!I�������+E,᠄��BU��*�S�y��w� aWWh�LٻW6���p��0�Et��O�YZc-s3sy�2F[^�BR��B��P��8�u^�WR�M�Gr�C>wjq�H9&�*�V`�K��er��O��hh������ׇέn�[�7	�^%��tf����j	ɧ[�k8��w#f���{�O� ��HM1���uCL��%��1q�B��)�\�U�*��?��j�y��wI%���LJ)�-�"%:����{�ͭ\�ɃP{m)��r��p�t���N��8�91���1�w[�Ҵ�̬t���(�~��$�?]φg��_Xť��`�<>� P�X��\ۋsݎ�N���傎�9 $��e���Ԇ��C��+,Ǜ�
���"\��i	X@��)�'������";�B;��0��F�K�.��nw'�����j�_��<q|�S:/N��� x���Z:m%s�ӓEVA<��1Q�W�/�B��10qq�� ��1��F�h����V�{*sx�	0��Խ&��\�� ��~������|U̍���gG���rݾ1_��O:��"�h,_�7=�׬��c�"�w�@�,�\�5kӮ�=�$�F�!i{�ȴX���Tu��Y/s� �		����ō	_ydĈ��Ջ1�Qf�sQH��GiW�k�K7֩0�a"=Np���4����O�I�s��fKO�����M� ������B�x�sV�/��9dq܍1��C�xDS  %�(-!:4}g]g~�!�C@�V.�	X4�(��g�W��f6�NJ������D��M�&*��ʉ����<{�]+�A��g���p��Y��63�_�w��	9p�<ѵ� GQ|�tn¸����cU���ű���?CO�6�f�F.��7,�[�ǁ�dO����.ol�^ĨTC�t��F.^�֨n�3/�E�N��7P#�"M��Q��|�P��W��V��vK�-��@��������ˉg���f�#d�6类��n:~7�X9*1�S���؀`0�ϩ�,k2��(=�]�}_�~G�}�;X��2��0$ ޖv��Ip-I���8Q[�=X牯MG�< ��j ��bp4c��ad��QpQ�։�b0��g����x�vǓfh/��QAS|:�ɾ��%�{5�<*xc���<�$��8��L_����,�]^�>�����g+���b�E�-^�ٕPŬ���aڅ�=��"b�&����C�1��De:��PЇ8��r�G3�n��x�GI�0�v��S6�� me�p��(�\���9ߏ�ԙqZ���NfWAHaz4��Wz��V ���yV�TG�jQk��}��0�g4)��o�OG�S�aI3ɑְ,�o�X�n#�G�T"V���ыiK	G� t�
�w��*Q>
�K���0V��M�^�j���S���� F�7񘰖��K�λ��ޓ΅#c��"�w�u��h���f��W%"�\Z�H�0��2��1� ._G��Gw1	I��\!X��;�,%�ZGeN�g����?�L
�<P��z����HJJ�@bN�8��l���j�~y�:�N��ɼQQ|M��4��٦���m�/j�.������d�Ȩ;��(rƂ���iʂJi�a��}�&�O�u8k���| �w�u�pJ����ƨ9T�T� �'�e!2`����Ծ�]��Ѐ���� �5��e�"XU��#J�ޗ�p��4VeظAN'ad��[��|M��SGH��tl>�o�a��t�����j��;������u�kπ%�|�*ub�&`�g���-{�Ok.�$���n��(wç��Lכ��'#�~�uz�6�嫤+5U��KC�sȭ��EC����o���w哵�5S���;sH{�'�F?_p�˺MB7�<a���M�#�ٹ�	t���~/%�Zʡ�4x@1�$,�k���M/�X�tWiH��zK	{'\q�	[3ՖˋP1Tc���^?�����E�Y���}�Bt)����r�{��/��*9a�t�S�L��
6"��l��b�Lԥ<�K�y&w�c���8��+3�o�qB�tw^�&f|P�ߚ�8�3���9W��*v;��<{�]B�8�HE�	Ǖ�ۧWS������ixՓ�K-#����Ƶt�_�n�����gʐ�l"[��A���(�a�4��fBc���亳NT���C0�Ԛ��O���0,��*l���)�i�ڠ'�z�S:��YZɉl�!fHBS���Y�G���zl�e��	���g7'[�e��m��#N7���JS��\H:=Ӌ����,K։05^x�	��M�t��������9�45��<���UzVI=Y@��]�}s���+YɹVY�َ5��cv�W�$vO4�%Vm8�}W��]yr9�N�r�q��R��\yu��ST&!~��o��������h�a���?Rb~�>q��Q�;gx��_�$��*�k� ���J�����˅�Ųp��x;��x�a���s�)��OOt!��<����8�ňs���N��;�gQ	�^�B�7Z�V=HNB$s
���	��E�Z��KdٳB����-k�p+]�ǎ�T0��_#3DU�1�t��L�$����G�ʖ�D���UT��>�r��mt�{a����i|�i�[�'���G�|ɒ�%�p)��<b ����n�^و�.�5p��e���+�bg8�!�ݴ�{\���MC�m�.�A����=����-&Ũ�d�����K�W�<���:����ƳW��H�a�����6������S��J���'�C�!�K�I�	M��^��&�+�o��1��Iq�e	&" �n�,isN���vM�06'5h)&KX�������5q� ��!��	�Z��H*�62Re��#5��m�.|g㺏1�C�TR�-'I��I�f;:�5�`�J��)�����r!C�<,3��m~�c�Gz4���224��Ϗ/\��Kѡĝ�Fw?�n�דT7+�E�)��j�Y����c�P kPZ?x�%D��v�Z�XX�U��?�	UA&Kl Ĝ�A,Ԍ���|Zŗ@t/�i�l�x쐳���;^��<<P�8��ѝK��~ ��΁I�0f�����Vg�v���EO�H�}������Nւ���W�5g��صv��	ܥ�r!���tk�Rp2�kHwHK�ڈ>M�O�n�(���b��bB�����N�AST��"`���?���n�C����wZw��eҹ-"��W`$y��
X��@����cΨA����������W���:QPRw�!nέ�k���d��y�K܊�c�]ߎ��Byk��D�c��W�Ţ�M����-n��e�e���ƒ�Kw� ���y�|�t[��C9������	��M��5��4�Qw���nfd�#�l]������m�
�P&�L>����e:7Z���>�a��3Mr{��UA\���9���W7w�U��Ս6�p5>i�݉�L�/���{Q�>Ŷ����aJ;W��!b��Σ_k�dඬ�Y�*�����`h�R�l7���y���5��'�.-ĉØR����k�k$��=ݴ�����2a��'������ql6�g�QoY,N��,��ܹ~�P˒�t��$�П�>�|�-��
�Z�& џ������ҭ�"y9��r@�Շ��;;J�a�fJZu�q�gr��:��R�G�SiS���%���-9��zە�I;������{X����}K���漢�Dх{���v�o��F��̚�����@&������� �_�=�e���m���1^��c-q�`y�BP�e�1��6�E�Ь�Q�"�aʵ�����m��U��>��0oq����O�x<i����+�炀�����n�У��ٴ�.uh�"k�_!��Z�b�c�+q�.�Hթ���C&rP�V}�Sm"n
��R���8̒ra�Δ��܌���������ߜF�	�z54�*�'�E���ZO�oxl eI*9r��u�2����tN �	�NW��r��XT�������كw� )xF
o��[�-�<���'�X888�y�RW�BOZ�U����$�q��ݐAf�x�^#���]8^J�C�1t����R-K��vS�Bh����<:�0�$����&H9�hd�������勖�X�'�%�/��?Nr�D7��m�9��8��.��6����Ǉ��H��
�j�Or =hdwz��串N�c�-����T���~�ן����Phe��������FF�+����<�pF�3�B���I`�Yh��"0 -���H���?YzL���ƾ/����O�Lg4=*�4
��Y8Z5�Y��a�Q�����٭��qis��s�G]l��z ��l�c��lt�%���:���@�nI��u�;8��&#A�������1qy|�y���4vo�z�T|#�#�GnoK�h��R����L�f����ꮕ �g'�7�F����n�7'ߛʌ_0%AID)˫NdOI7��S������4����v,���dY0ކt�����ݍ�!����>,j�d�+��>�^�Q!N�H-]��b}�/-�hŃo~�r<���/�'=�(�5܏��̊��� 0H�e=T�|靘��3����)�(}��߬yH�X��D��7�磅}���i��	]d����,��4t�L��VU�u��6�ܲWc�]eʚmBW�s1@��|`�q�	�^�s�7�z��4��_�$�=*�_�%�T�*P��s����WM*1�>�O���rJ�K�T�����פ����.��ðX8܋V������� m���TW&�VZ�Nގ�d�4V�#}�y@R<�eҥ1p�`5c{c+�J�A�j��S�{Z����F�a)j��9���Iţ�J<�!��A����z��~=Y�E�:	�V���x��-d�	3�zQA��L�X�ҥ�k���Wt����uX��Q���(y	���e�]�Bqm�S�DwV'��$����h<���瓉�$v5���"E�~Jw��[�ƛ��Yv4��˭ԥ�x���[�w�J�\Y���{+�����bZ���w�?�L��H�q����2e��i�Xš�L��lH��j��^{A䆟Mjۀ�����tp�"[�4������D�E���a{�>�/���R:�l򀮆��Ɇ-�NK�m���Y]xj0�����gZ)����0�}u��a�,A��\Ϸ�_���Q:�kF����(�#V��B���B�(�z��ԣ��Ѓ�M�,�N�tT,6k�5�_�T
?7���>8Wj�3�WJ5�f���0���m�Q�o�Q�
1���x����OUL���;����+��4	\,�4�G���Ԋ�M���['B�ј�G�������7Q{����J*lwtK���P���톀:`<��n�"
z�C9�m-�vu��$����9o���7TT�y�����8g�����eh���,�X�[߬*�'uA.�9�)�_{��F����Qyyv����@����@�Il�M�n_
�"'����{
GD�����B|1L�*�W����Dǎ�k)�#��Q�J����<b�_O�Z�����q>|�w�k5EW�G���[*��t ����p�,��m3=��� B��Vz�fHX<J�$���nث4���:<)��G��j��(�j\�^�Ft��N��V�#�H�ѧ�[a�<%k� x�a�6��%?���da��R
E�.'~ݴ����vg�v����D�˅�z;�<t8t�˽�7Z[�`m��WG���Fy��t�D��>�O�Ie	�x��t�y8�6#=�,S���w걇&};�|ߠ�ɍC�a3��	Ƙ͟��I�� �׼hi�"4��DY?���xk��pY+O�SP�D�}�B'�4s�^?��^f�7ۥ��$����e�TE�������K�>�eM|�;��>	���p�+�Q?��v��hZ^����u?�4�j�������m`{P(c��Q��B�Z
�2���秶b�"���L��:/!Z֌uS��������T�
S�d����7+n���7��xHhfoh��I]����IU�ѝ�-*��#���FHG�[�M6����JF�+��>�0�ݥ�J�;��Nt�	1�&*谍�B݇�i8z���*�cU��X��n.�V��%-��EsbQ�"�(�d����aU�Q&�m��ZZ��l>[��$�����D����>aC=��"a��*7��E��r�H�d�o�J�o7�rk���`�f��ȕ��J"�ϛ��5�� �YA3h�"��Q�j���T<D�X>�u�@��@ X�h�/yj�(�%��aK�#�dcoC�C��|Gˍ@}�%͠a�
����`�g?�zȥ uH�^*��L���,6�0����<�k��r0���V���{������1������܇��Af�ْ��
Ҥ���[Ȇl^�ٝ2�]�r�0�?)B<�RCm ���dx�	�k�E��CI�!/�d�x�ZasP�y^Q]���P��T�웑���B��f�\��y��"s������F�=��Qb@#`f>��7Ќ3
h^��+7�T�x� aP)���S6	�h&P���B��;�9Eo��:�qq���� K�-]�B�����b�Z�X�	Z7��Zʐ�&3��"������/���b��.�RM�Փ�nez�W��h:�������`�0��<'-��3P�/���}%�>o�c�\ �w�ۿ��|D��6-ڪw�����v.7�g�T�+c�Nx �p\�ݳ�4] 5�f�@> �=�=z%�OQ�ԒxbT���k/�rn=�%+Xɢ�-�?W`���� �~�{�˸U+�{{ߕ�V������BϚi�~����ƶ��Mv��;�}3�v79�q���=$�]4b���w�5]��ŁU~���;��b�y|D�����t4����ݛ?��Gpr��8�uE�ok6��f�D�-⽝����L��6r>ٝP[+L����J��zN���qH��L���t���-��kq��!���K���U��9�0�����\�cNK�M�m���,���'�����Ku��mM�$=����1����,�������\^ˆ~d�tѧ����sYwr�BNXA��`���b�$n�Ğ2#�I��C�\�ʑVO�
�yH��H����_�"`7�.6�.�l����tD
���"�<�������_2������������1��L��5<������@�)I1��܋����c���5��fx�e�`���^7m{;\�~�f��{�ww>F?�\�%����"J��I���#S0���R��nX>j��|�{��o�	��y1s��s~��9'�%�)t����0�8���g�F�/���B�9-=�Ol�8~�l��"6��Nغ�����0@ӥ5�/�������8Ft,��E�H�8AE#Ӝ�0M�9�){t�O��J�d�^DD���j,-��V3��Z|�ԑ`�s�z�c3;[x�����xb:���'�A6�Ŝ�1��5��_Z<��:��*8Q�2�$>`)�]A�A��\
�������s��#����<@k!:�F'�];KY����x$��N�=/Z֪5ls���$�_�Ϙ�����ũŗ�F..y�\��@�ћ+�!G~<���~�a&�0)�+�޹�U��'��U�,e/iv"��m
\,���S6*�d��x��������j�]?6� >_�� H���t�ĕ��!<�WP{��䴺�,g�V	����RPpD���m�����vD4��u{�'�}3�/��R����: �) ��	���T��bv�[3G6=Ԩm�fx��B23���Ϛ�b��ݮ�P �՗/
i8	〜����T�?p��W+(�����b��v%�/�p���j&���d�M~�/�=���Xby�ݑ�i5���E?%�"<���oR���{�V-�r��q���a�n�{�!�+��]!�����&#o����Tf�È��?�EC���_��u����#��Ĺ���Y�"�"����4�C�+��=9#��6��<�u�9�'Puz�8�Q}�l�g��ߏ���E��&���n�v�
��QU�$_��I��a��&q�����6���O	A��r�����!�̨xq\`I؍0QNZ����P�;��I�m,9�(��1ē�'h�<�ֿ%�MA\I,�2C+j�1]�n��ܸѹ�r�:�:.�,sSL}�6i�x�v09�	G�^MzW[��K�*� t���)c}r�3���N�י2������	���Ի��y5�r��yɿ��L^��qyf�������&P%
@w5n�"���9���7�h��x�/�^r�m��$���~����o�m�׫�UY@7��;�.��$��B���)?TԘ���P>C��f��6�#�&��fI�1�c!%cx�G!�*�{��1��V��DK��po�e�b	�I�kyb�����Z'>:2~(˖��W ��E��WQ���M���o��u舦���bA��q-U�RD!p봅��+�t��R���'vX�иň��a	2�T��C���CWEd���a�_F�N�`���#W�L�)���l'����K�y6�v����I���X�Wh��u�]�.��I��O�9>I�[���RB8^���+�z�����q�y/��b��ß����pژ·4�w��1�w|��ӯSj���0opp��C��׬�&�.x}�� O�<$��)��P��Ϳ�F��4zƗ[��A�>v�X�i�c�"[��D��;�_�9R�ō{Z��a�e�UK������H۹�
�'jOB���k��p��5̇�a�L�Û��%�b��zPTq�#:�ZG����}G:�a�A}a�!c�;��CL+��;�h�G#&T\��@���D��s��u���A�
O�s9f��<�����E_&ca ��c:ה��?�!��~�AA�m�%��r���G��On��"=5��th��$���`)_��(��Ƈt)�p���`����`���K{��(=&�sT�?�eb�P'�ξS�n2�v��³3c���֜�36���)�vbd��23�p��3'����)5�+
ə}}3��'�غ���i����'��2+��	*ྉ�
m�����g���[a�lH�v����Jd��X�7k��Yl�#a����TV/r�#�zw�Fl��m���煊1���JR?�d�
����.����.H���f͌�-���,�`" �$�[,��q�G��9��-:�P3�y,�ܚ����>W-��Z�C��K�&�2R�,F�KYpSG��4�ߞ��-jQ��E���H?K幊7�rn�Et����'��z�h�s���v����K��ĝ��V9�￴������;��蹔�R�&��<j�˺� *�0mj�%]������R�;�T�ƿ��5�;�>�`� �y������*ۈ�/��'x
���!P�HU��J9����HĽ��\o@�L{�r����]��o�^�sG��ks[i8%�(΂����քbV&�/������!eG�X�E��/�UwHNM�UFR���]5&��?��M�o?M��sr$�<>楺(�-Q�j�>4�5��c�̭|���'��h��6��|�ANT�%�f�����\o��Ϻuy;�a��p.��:AJR��$�V9neūXȘT&R��N|B���	����-�ط�u���xX_��q��V�UZh�+�Xs��m��E��h���ɛ2h�o�%�P���!����9��+5R]6<U��5��n����=�OE�kL��:D���<�Pgʆ����v��
��?���s=CCk��(�q��T�= ���/�J��loݹ��̻W��x��Cʔ���z`Y-��o^��*���Ԅ���F�P� DU�d��.kb5w��^T7��Y�-��md�#���&�+�s[=T߸��l��$����*ќ䃁l'��S)^�C�CC������r�gTA�oq��Ɨ���	�&��R�_�<�+D|@	?}���=	��U���_?�� �`L��q���� Y���k]%���G�o��a�v�p�B�kݶ0n�;��o_��Zq�����%��x2�����y8�����ͮ�F���rzϰ�EEO��Kb5/�T�g�fN��m�O38���04(���^��ѝ�rFB�,�������WЍzߕŇ�rm=wQ ���K�T�m^8"Q�z��m��hDw�ᰉ���ܭ ���7�[��l0�� 4y�5��fn���:ٗB&��x�~W�&�p�+��)ҸeuB����B����a.�M�
��`�D�$�7D�ϕٹ����=��$�'q��[��N%�Mx^,��f�O�4��Ш�U���s�AV��&{�R9��,�g!���b��%���{�5�y\��Bo~��-ϝ������6m����f�p�o+(ʄ��-i�+�R1)�1�:��ڞF)iѤIㅖ����§��)�'m���`��2j��j���Z��I>��+��֐���!��b�	"��bN�KM$��P�\�,���G����.g��V�[��;c�Ӎx���0� 6���z�( yZc?��l�����I��{��(:I���:��P4U���oO������c��}1+,�W'x����)�X��S>��l���'׽�=d[`�r�e�L�),��.�It�W �j�H�_.��;���|,�64~�3��~N�D"տ�5���֧�[<��0�w��Ð
S��sS�t`T���V�&�(��9'�� P��R�@�-�N+']J���o)����i%�Y���κ�������+��KRaV��Uߝ�
^�ۮ��_��;�"�t��qv�qr+�`��8]c'���1`��)��q������JW~��OxY��?B�/g%��YS�,׋�3�OX��,�D9�M������*���3l�BcÞ�G.@{M�����Ђ��;�S?�ގs�A����K�+|��h�_���~ǝH�P��YW��U�0����|�[H�Ԕ��+��Ҕ��"��'��ur�ED�:Jh*xW8��E<�<�r��bEm�@{WQ�ũI܁n��Ou_@���F�dqt�2B�{�=�,x8�!���u~Oo� QT�In>$&�q�*�qC��0��F@�z���t��I;W��z�m��������C������8e�6�GK;����6ޜUn�Ny�B��}���c�����V�����0~aX��9�%�P1�q�h����]������1�B]%�A���|�i��gX�<�.�"�tfg<�/�؋|����=��;VW�d���?|�c��@�^�nA��s�'8���7���X��sH�෬P`����9-�J��ӹ�FoW�y=ՙ���'W�mb�XA*�J�U��[/G��ʸ I���9�Ez
��N�^[f�&��di��۴���$C�Ɣ���܌δ��i��]j�����i�V�VE���/b[�,P�
�R��2��kN��6�ߏ��pט[%F�'䰋G#j�U:��wV�n��� ��XK�18G9ԩ�L����
<�����s�kjKPp�)��)�wh�}�7q
�>MiS�Y=���V?���S�����@5V|Fi*�R)[�}#�б��+�F!�\�c" ��΂*�qklJ���tC�l��n����.��N>
(��R구l���\Ĉ��ZC����SvA�Zܷ�aR&��ߖ�Zp	�F����JF��p�UH�|e9k$�Qƍȼ#4����4��q�&��͐<���u.0�[M�EjA���%HdE�e��G�]�!�]�X�48r�X��O�_���3�l�j2� O���r�>�ԝ�*$UO3�_ɾ�����k��4�X�N�f�b"��4`���[�C/x���?���:��4$'с�QZ���*3��g,P�����m^
��)Bб����e�J�ɑt�k���f��G承��\. ��e��F�O�_p��+��s��,���
́t�S��� .ii~m��ܱ| � @�M���k ǖ\��lb��8Q�前���ޱj(8a�q��ьF�l2�2�py��� g��V�Ⱥ����K�k��S��!���S�B��,ǲ�_:Ǯ�6�*�6G�r֔�]V���K�c�������8شQ�3�e�`���F0�_�?��J�+3����zm������!~��4Ĭ;��W�E3ZӀQ�f�<�]���Aѻ��%�7�.N���'�y�W��G��F�ʍ�C��a`}��]$���X'�u&�`��m��N�+�ʳX��跾���A�Ǆ������x��'S>��/�R������qak��ɢ>.�w�C������$Z(����$��.ܦ�e�
�5q8?���$��w���W�ay�4�tG?���uP?,��q�^����o��.ѳ�.*�E?֮i��K���,����!�K$�Nl�������tVZ_��@ĕq��K����I ���j���	���If�}B��5�r��ժ�{���?qK�}�s?4e���#�E���\���T�a8!a7�|cN<DT�,
zX.�h�k����f%�`W��T#3M����^MAˉ�#$�=�rUK-a9���tW���RV
P#�6��۾0�]jx\�q7ح��>�EW4ǩ����9��h!t�!P�.��j��/���,9�7%O�$k��K
9�ý	�i�*��t�/�!���t��/��S��΃�����o����Ez^��e�"��M��cs=F$	�
�>���FԽn��-	����Im �o�Oti]u��	��t���f���\8����H��4��%7ݞӎ:wf��9a�'� 0+�<�f=�BE����(N�0�ȥ�����ɶuou|鮶6੊VA*o�'��鮱����t'ꁼI2�K�����ϋ���!p�\k ��j�äZ͹��}�G"��k�^G�c�(���i(0,S��ap�ā�Z���Ƀ2h�i4)����hS�0�=ųor�LV�湿jB�S���vh�~NN}+���y��Q�N�D�Q��]>l�����؈�1v�*W񾛢)��W��Ģ$
̦��>2��|)���v�kP���d%>YՏ�J�HК�nz<��ú�{0����N�w�6`?�A��^$kE�
9��~^��@�E�P�X��#[W�!s����s�����ґN����9o��5��/>�U7z	t�r�0Dc�}~�����䰝�,Md>��u���Bi�r�4C(���ӢQ���� �q���%�r/s��?d��O!�
A ���z$�DP��'�w��F���1�ӗ3�B�m�ר|Z׶W�@�W�ğl�&��Y.���s%0BT�3K���m�E��I3�J~uف"M�O��n����y<���-�AܨV3l�cơt2�HF�P�޵��f.�$B����p��_vj7Yy��]uû��N�2=���Kp�W'3��p�"h�G�����I���uQ���h�u���ç]���_Ż�sޔ��Y����hJ	L2@��nwyC��޳YOG��O����!�t���#o9"�!�B�}�;��2n�B@(t�@T��ym@���Ї[W������"ϣ��UGY;�^����~�obneM#���n��d���[��cn�PІ��w\�R0��c闣[A#vc��:�
Z���%�5��D����!��p�����,n��A�E�ן�OI 8�Q�w��'Tx�j2�:�oSD��:tz�]� O��m��/-0 ���4cPr)E���*�ԳV(�Q�6�d��NF+�j���eӦݵ=fS�H���'��O�g�����~�Q@pOv��?M�m�av��m��~�nPWB�Q��!
�F�v�y�ב������*w�$���I`�s~9<��;@�l�ƫi�e��&��)>Rg�[�5
��\����� O�n )�@�;w鄾��zPW>�n[˖G�Q��C,Յ��'%��y�3Mn�I�����jPM���\��`�^�a�Ľ�I`e]9p����d�8!�����Wo����+D-���E{SYB��POV���v���­�O9%��/���L���F��Q�ä�Z�%	K�� ��K��K,�ҵMf��
9f����Y'�o~GL2	��'����)k݆�r��'��u���O�b3N3��N?Ӑ�嗂=c���� �j����xҒ�m�����ӅU����|#��v%�r]�8�(�E��~��E��zn�$���@0vA�:߲��yIi@�n�r��4M7o��෧�aXi��Y0 +&���UW=���D{��>O�*�\6jY�9�fhv�e�{Gʕd}�j�n��v�vp�S�$â�����c�uqX�,�U)|]�_��ՓFfM�4��&�.}�� Wʇ��h'�%h�����0�J!κ��"�	xq�*��v�&x�Q8����������i	�*ݵ�(����?%ʚw�-��#�Q��#����ӣ��5eG��r#�[�(�]��F�����:+��"�
�(0a���]6Y��e`�5m�UbX^G)M:s~�4]Ug]�`���b�<�����
��=������X��_�.��.��W$3���R�-%� ��{���j����^Y����<��f�f��9d�W����R��E��HC{X�/�8B�y�.��!O����39�D+H��_�!�ﺟnnK*pK��W��r�?��4M+�eѳ�z��u��$9���:�~h�5J��о ����m:o*�, ��SڨIQwf����:e�F¡P���cT�5G�L�ü ���j���]��|̆��E ;���puǁ ��b��V�j�G�_�k������?Y�1̹�s۰�L��;w�M�ω��j!�w����Y7QQ�sa�j��S	�Gxڻ�,V�y-�H�K'���7.~�RZ�c�%���<xB���i'霖#�4O�ܜ��E�׋�wemS�N�����Q��@�?�Mk'�T�ߌw�+��p�j:-Q1����P�K~�L9Z��6	O��S R"r���tl~ܯ�������g�sQ�)���	~Ѱh�#V*�V_��>���W�|�@�a�f��D�cݗ�������G�:c'��)���)�౰}ٶ�"�6Tq.��.0�J���S\Y�CC������KX�7ח�dS�6����*���xu����[�P߲���_I^}qBU".�!x��ܐaZk���T������[l��9�닾����Y���|���<��KG�
6��9|��:�����Tf$A,���h$����������>���D�-���XQ ���2���p��^�ŪY�_1�A��Jsxi3'���#ڗjIC���+�����쑮�)��e�~a���������,��XB����]�W��w���7k���L�P>�h�)��O�c�r�ky��cV"}�2�xo/j�����>%a#�Iv�ϙ��Eu�k��̧KEr�6�d�V�٧�;��������I���U�[�����Z��T�Ƨzrͳl=q`_�,�;x�OU�*��@�kmfG�L�i����]6��t�a/6(ȑ�n�ґP�1ڔ��A��X���ͤ�r�-���K��i�2�튀h�9dſ��9���W�	pW��t�=ě�%�]h�S���<��-nri�� �/��b���F9a^D����_o�0��(�����wƋ Klb#�L�� �)��'���+����F�! cDN�����#����z��������!�g%DIA�۬��涱*���B����D������ �I�B|>N3�s!��a S��dlj}���ë^=Q��8��I}N��h�:��(u�j��+Q�E�Hݾ��ɥ�V��}�z)8���:a�!x�p���R�ild��O���6ޜ�ue��t��F�({fr&?-�x���6�ۭ+|
�����>98<W!���Κ�Cj%��ïq��g�(��wS�* F�:6e�s�<�>��*g�P�\NȟP�=l5�G�L��|Ù���h~��� Ăǰ�@���e, <��^HeB�A������0a�#��mr��vL�W~.��M���k���w_� +�k�(�N�)���;��i��TF\�����sLDy%b2�u��"��b���Z5t	���+;&���6�.`n:�_$�/�[DV�{:���!����]H*z�;�@P@ߗt�Ri&�{D��~݉R=�>)�^*з_]�`�a����?�����ЮXZ��hTvrX5�p5��6J�tl��O��G�S�r%���"�ڳ`Ng�p��O��8���I��(�r�5G,���R����uמ�+���hn,���TDvİ��,�Qf�G��JG�����r�8�S����#�+f)����[�����׎�av�K4�\��XM���|��QF��&.]+�A ��&�?<�ĊP��Gj�����^�VS48΂�.����Iұ_��:����n���1Z��e�[�s���Jna�i�g��,�Q��=�p��ǰ��g�Zj6�u_�e�!5:WE��bw�&îԚ�m�B'�C�a%�1�1$ѐ{��gw��i`�-N�8�mfU��P��-��7"�u���on��y�I�4�j捁J�Lmh̆��N� ��M�`��Qu)�ļr�]7��g;b�{��o��>���Xd&@-YګJߙ�.	D��	��p�[ڭ�j{�p���Z?q(o+M� �߽=F@�Ai�n��^d<P��c\�������י^a<1�������#0���"��(z:��Ȇ����ש�������=u5���ur�%%��"�-tJ���Zƾ.� ���-Y�R�9��*r@�	�8s�;P,2�>Wdݵ�KV�}P� ��)f4O�8�"$�����9�FEr���ʓ�)BhT��IP%�k��h�6��d\`��I���V�Z�r�g�X
j���#�F��xE� �r�5�:�~�+m{�?;�
vN��R��}��j�-�0�_������c8��<!���u�(Ef�_w��n1|�l�����ڋ�X�V�u� ��"4W5m�P����Z���Ll��ˠ���W���L�_7�u ���/S�"�8Q�:۵t�9���f�-�q�%�VW\�Ú7�%�.�KD���od?Nsk}�����J��1�2)�m1?��{����3�y�z�������H����V�Qa>�瘤����� �9
�c9���k�C�.�p��|�v�"f�� �zX��)z��)�F�,����̣kk�E��^i�j�vd�%�u���]i�WM��a^v��$O� x�����Y)zO�f��_���I1�(?T$�N~?{����`���kh2yb?��8�/rĂ�0�RT�v��!���n�r�(;?v����7C��uuƗ�M�#z�� �
`Rg�;B��e����L���GQ�����E,���˜�"�:����NQe�)����)&����t�}�@��~�8z��T�*,<��$VC��T�FF&�X�;q(h*N��0� ��Ҩ%��{B�Z0R���d����i]E���&���>Zc5?6��i!K���]���>��>�bI��#���a���}۵���ޙ�в�d(��\��&���i}�;Z�Ӡ�w����U��?Y?���s�^��aԜ����i�&&2QT75��j�#q]�˅��׳L�_����X�rg��*G���㥼L��eaq�n�ͪ�P�ߌ0�4�;�S�	4��o-B�.ķ���W���W�7rź�r�t�ƻ{��Y���́L��@x�>��^����@ ��YƙU{'Zg:�_G.����j4����`��y{5���@E3���k&nȖ��#��-1�՟2be�q-��p��5�>ϑ�K�����s�(�!��Co�$�>)���_`��s�E��J�ń� ��IH�iͱ�d��IL~QY�{ n��$��p������}f\qn�H���[�2q���S^��E�}������Sn=֐�kC�߲��<j�y�0�Z���}T���?�)�ř�7�B.#1>��Z��|�%f'#	&& ��az4����O#PM��o��ɓ1Vm�[fx�ﲧ��m�sLԾ��pWzH�i�L�m���s�F4��f�W���˖4W�5��"j���ð �1.���1���}V��Ƞ�Z���:��.\ ���ϱ�>GHb[s$�A��Q�k�SWt�HT����@8����Ά �����b} 헯��E��zDP����0����{.���l#v�?�#л� ���G����l�T�x��o�����L+�:���y�_����upp!+7f��q�5�o�e�/J�ʲ�bYٿ�E^�n�a���4@
@� ���팄�e�D3nz��^�����L�%�ɽ~r�Tn�6C��N��[�hkG�3a��Sl�sd���"�YU�W��3���V��"̌B5h�<C���iT�{�ʶ�isxE��g��.��P#1^M�[ol[�I7������=B_���+V!N�l���s<��i`�����&s��{�xdE�^y~m�0GW��(�7�F��3�A�4M5��P���W���|���]��7MDV����a�V�ߘ���YxO�GB*�2ό��#�
8�S���?�>Л�6vU��Q�T�R��[G��Z,W��M���N����|l�:t�bйC�t�| �S�2��g�ì�e�}\<~@�
g�;�6�h,�q�v, �k���k�����T���ά�W�8���y�uM��YU}��0�+.�<3�.t�F��!�aY*�s6��P�~�r]�]���m�VX�u\���4��0�r4���i�o4��9��X�*$�S�`���)��`f{�W�9�"��E�,W��U�� �S�7�D�E��ʔk�#5�\a.�('���A�T�|Q,o�bP�TQ����a���Y�*w��On_U㦨9�8(��F�wD�}�S����WS5q��Py3i���"���*q��!M��l��"n���L�P3��� ����ݩQ����z��Z=.�#�ϡd)#'����>��@�e���-����A�nʔ�th�c�cX�"�����$�S�gkv���e9q�	.1������ u.dj��և>e�� {*��j�N��p�+7�l��k#&\���#߽;��7�*v�eKQ~�]�9c�����b��wf��b��	��ݜ�W�,k=�ǰ����W�m��_�B�v'|��S�*M+�r��Ȩ�rElE�H{�?w&�}m
�9�g\P]+�i܏0O` blZ���I,x�\-���^ߞI�����j7ى��>۟q�.]I]bn��.I2�j�ゆKAi��؟�4�j� q�sV	�T@�����I���w�a�E��a]D�%0����;���}	�r�(�L��6Mw�SĹ57?ݖb���踚M �M�,���8�]ϰ�8iѯ�p�̉�M�C|uןMspW����F>�^g����a��ǏUU�;�|Lhb� ��z{�2�(�I=rz{b�J�g��zB�8��p{�v��	nz�ۘ���V�=M<-6+� "��_��qG��=.��H{H�?w/�wJ��G4S���x�����q�L#n�f/�p��GpcT��t�g��$�� ��)�̍��r���9є?C����^���W�Q2����2~V�S�>?�^���vm��7;I�����ͫ���I��S��c�Ə��hng���_�Čf�#ۃ�
�{P��4�m����Jwo�i8�|�Š�%ޓ�'t�g������t=��*��!3��^eߡ%;eU����Uȁ��A�i	b/��ff��\���m��d0�tOv΀-b��T�z��h(<����f�ᾘ��4*�Y� : h�«[�|1�^�S8�u��P��Ӛ_w�Z�ʓ�bo�ł���/Q2��n-F�4��s1�ʢ� �C��P�rS�K��q���<�	9�����6EyQ�Lֺ"A\�\��G��-[LO���[j���ۋD�A,����^�u1�yvx��� ����E��c����T}Iĉ-�1jC;��BU����rqvO�S����C3�P���_��R�:	L��t�(�+t]S�K������<P�쩂Y��ܨ%������k Vj�2Z%�j��
7t�l=�{�1Φ7�VX��Ӱ�f�����ŌfO���˷F�iJ�;����ʜ\��l��'?����JX1
F S��p	?ڿ6�7��q�)�5�r���d�d�tN/}�OTim�_ �����2��.'v4��?�cf_�U���Ӈ'uhٚP+)
(�d ���I���c�1����i8��D���7��s �����1����<�����f�u(Y�Xc��sWp"�vp���'��D.�<p|��������-�:�$����C�b�C8�)(��h�|� �ֶ86�F�IC�Q�ft�0��һ��6RJ��u�c�p3:��E��N�5ƍ'� �
�sZUN�۱x�����:X���Xbq���)N#�ޯp�Kb	�S�|!"��P6B}=�M��h}C9j��O��
�ԫ�8K-�7��v/� D�} �{�{��.� ���4���'���kr퇭�¹t����Q���sIR&�a|�/`�@i afx�����)�7>�0�n�K����]�V����
'>�NO�5:4�}��F�o�[����`1D�++�pp$x
�%��ه�k�Y��3�nj�&�A{l���w��5�wS���1��%fO(Q��N�C}P���Y �B�_[�j�������I������dw)�冀�aN��{y|���Sd�n���T!["
���%5-C#���X	rt%�2���a��&�REc��p;tg�Kp�vwɇU������<���d+ Ox/�1��/%��mn�xR�\�	0y�{S����lT��Y�ǰ�5���?�N�4$Z�7�ػ���3h3唨��n��Xkz�,Z����8�@��z�*���#t�M�kvV�u��$��\X%��H�͊C�I���(G�`��Nr����?�ۘ.At���JluQ%�5�2�e~��b=1��6[�:���#�v�D�4{S��S$�.WGz��c�(B�U�ܬ��\���&��W����✏��k$�v�y�I7YE�iuٺ���"���K��0z�$��N9��+� �~�V��ߡm���������
�y�<����<��`eJ���P���~IjS����R��e&�)'�%׵�������|n3l"�w��.���������xk�$��lMh��$��,�u@�Շ�>Сg����4UV�M�ՀB>:�%���Jj�B�o�:
����lF���&��C!�\�X�k�O��V8�4'���&M��ܾ�0�0]-�))̾��$HO�p���v:��� �~�����ߜZU�df��z�8���`�z5߉������}e��p��r3�����t>sgYQ=��.d�-ST��ךM"�(W����4����H:�trO�"��0\����@�$A�{��d�J�����Z�dQJ%�~�Ɠ��!��FMa�$�B���p��%ܟ�50Ms�Vq�6f�?9����X߳|u*�U:����Z}5}h`FWi\��El>7k��;u*!l�Q��[2��#E{?N�����\X$�7镬ggg�P��.j�����6x����bL'�I��u` �� ��Evʁ�4�.��-��;�!�Le&�l{�B03��g��� 8��	 �����$R��?1Xf.=}>����U� �6K�">�.CA��}ӷč�2%i�d��^Js��߱�m1+�����������˅��$�II�o���� k�5ª)�Qk��9?x1k�|�Z7V���Ń�ݔ����h����!��g���>�s�z���n)x�Ry}��\@�
r'w6*1�<�4Nw���R'��͍� jx�%$���`5�'f�-�Uoh9�����'�s��1�Q��<e�p�U�({w����3�N�-�l�9N��_�Y�0�7f�p��?���w;*�/��ą�����{��Gj�p�JG|9�6��ϳ���Zw�c����1,�s��d+��d/n6`��"��{�7�:l��sf$`�Q�D5��W��!1�e��<[���($���dM�2��V�"0����=���Z���M8E��}?ɑآ�9�g:cY9���fF�-�S�+|���X�j��������jbidn�i��L^��V�O",@�C�ڹ���6 ��ku�`�y�'�4ᅇt�}� "	R���^�?�A�6���E�s��``�qzD"(>}7]H���(� ЍF̊V�}r��e�$k�$�gCy6j9Y׈�jG���Kwߊ׀Թ�2ql`�:a�ѐ0�c��tX���q�jѺ��p�3�;!uј�$��U�N-���?[��ق�<��qu<�J������	_�8`c4��Ya��%y��R#��-ۼ�x�e���g�r�
&�$(�е��~N$e��=�H�	/!��+�D��W���]��=p.h~J0����3p�QK�R���H�8�Z豔o|��|�G[T�2Lʠ`�l��lu���)B@+[�������H+F0D�(x��o�0VY�	�����m1���@���1Bf'��W *	Q 'Z��kĂ"����"�G�-?	B��&���Ѱ�Oa�[��=K8"��?��j�C'uK{�'g�L��!I���>�&W�EB*Ń�MwQ���YRE�6l�\
dz���d��V�ڹ�V�!VZ��.�wG��(���}�XZ��Uv8�s�㿕��{g:5�J/���c�ja5�������0�\��D^h�m��S�k�K�ۂ9��Rvy�myJ�Q�YS0�4h�.KS��^��gm�:��hXRe��Gܕ1�1��╒/b�h"�_��.�} ���-�Z���Rm�M�iUؿ +,񗈬F�,|��<�#��6Y�QU�QL>��Ş��ȍ�%�Ye�+���pKR�|νQ8	R3P9��/�d�$�MZX1	�HŜ�d�@�ψB����M~���{`ƶ������K@(?>_�6ء7��S�MM����5�(-���(�N,��N��m�+�!�O�mQ:��������OȪ��W$�~�m�	Ը)����2�)�o�\
ɤ��`9R�����u��!�uѿ���qg�yN�gg�,��,)��t�d�vE>O��@x�p�b(z�����o�;D�"v.ve�q���cdYUZv3NC���T�5|q3F�ŭ夛���I�l�1{g�B�0��[��|���N�v��h;>�Ž	���m�	^<0��fI��d�(���TK�!��\�oy��oUn��T���b5��SgH�C�q&L)�w���r7��L��Y�V�)nEu��|���C^C��a���s�=k�.�����E}��䙻���nޥ-����#�.���ۙ����7PǍ���%��bD�������o>�i�/WĄׂ~�C�D�$�6�i
�/�kHY�>����
�/9��XOI,�S!ZA�
��מ�%��yZ7t�B�8����ܾ�)�����#�!�#_N%Jz���"7[d{~mlʦ�V�8/�@$�g�S;(�0�x���o�F���w��o*+���w��$#Q�@ _���!�~T�fϵ<cV_?\?��[���ǴgB��Q��,ش%�L��u�v��Jw�6L�;{w��5TX$v[;/hȞF���?G+4ܸn�O�Ω�L��N'z�p�K��r�ޮ�]VVͭ!������o�����;B�"��F�$���/ԏӟ�i$�`�-��H���^Mn�3�8]�ƒ5�h����ҧ�M-�ď�i�i��J+Ԡ�c��+�i���U-�J�A���5u$(ĉ�Վ�hDq�x������������ϱ����B��i�����Ӈ�+�J���f��EG��|���=>� ���UB}�	y�z�m�>q�B�S�%�tae�.jb�?ګ?���Tͻ��������1$��f�byC���ԛ����f�y�ք��^�D
4OzV��S;7�C��.���H�ɘz[uC��R\�8/\zb�W=��@Tl��2��۱���U|�>��t���,X���R�i ��������XG��Gf#aP���~�i���W�@�a!2:Cy�}��&	j��>h����@=g���'�g/��v%�2* �ߺ�I�(���Gq�%�8���SV!ȟ.'I(���>��,z/Y%���"��9�Hm��V���a��ـ};���>O���?dr�D�k�eWa��歮�Rv����^��tJ9���ew<�s�5�i'k]��.��ǌ7��(<w}ʨ6/�Pv9�'���ӂ����x�~�fl�9�\�S��u�(V��M��X��/�pt
2�9��U��'��uT$�	�d�xE���5�))�B��`��U���й��6������*ݓ�H�z��u���T�{d����[��<���:��!��KJ�Vb|~��ĤR~���������o�p����^)�nDyp:d-��G5Z�9*��_��j#�%@͋���3 ��}�����ʨ0e�;�jÓ|��ӌ�`�h��R��?7(�p�;���K��m�>C����]1�	��#���0Iad<8$>�Dr,G; uT�����☨��(-+/�����5��+!Bgl_n3�7�(:��#��>W��������!���z^�^䄗���ع�������nυ���[�s�ui�\�%䧪�옟5��H���e^Jv�vaڍ�@z�Jv뢀b:��3�cyk瀭��e����[�I�0��I����
v�V�+��	s'�����*eО���36�4�B�MQ�h%��7��_��U�n�����:(T���"{�ڒ�|(I������E.���NdPb���ߊy�?٪FI�.�	�xj/�����j:ޖNs����
2{���Cmĥt�z#��i�LA���i?���7~)dx>y�k�Tu�c��JkZq�"�< 	J.o�KO�1pz��cq�*���%���ߝ���<��G^4�����gˁ�F�_�?r̙��2�F0*�M�E.]CN���03��$F	�J!��Vѽ3V:b�K $ˣf&��7��9�ҍ�7��啟�+�&�H/1J�?=:�&�� JRhoO;�Κ�����G[!��T�
�J�C:p+����o���ȷ�X�@�k�u*���I+��s��L�N�b�]�w�PP8����-yL �QH	�{(Q̴�?Q����]$߉!"�v��~��5@np\>�e{��}Ƙ$��8lF%
GM�3=H�A-%@��p�����(I1�_Q�`��g!�nh*Z�,dw;b��o��-s�.P�k��P�g���S���=�8?�9O�7����n�=�lp J��$�}���~!�i�<oz�����Qk�ꙣ׋���������]u�xa<�4�Q`o�_<	������˙e�D�����$^<��k�ev1_7痓Q�.��a�H�m���`M����#�<|��,nh��}����)8�w��q��m���NH�]��b�`����Ay��@U(��U�n�p�DO�p{Ѻ�-���h7�̠[N����h��D z�te�F�Ј��~a��0��֧%�敡�?%r��4���c_/� r��e��r�X"�Y�nf׽��Hꮯ5���O�o��e�mǄt��s>
X�ЉdQ�ЦO��g:�N�n�~���\�l����d����V:����P�
�����"�(AM#�E�#��)�mSc�
�c1�~�����4�,.�Y��eE�N#j�A�v�hJ��@l$��c>���cn+�WJ��CJ�5͍Wj��4�nX��j�
a=�h��;����Oլ1��*�:�4�(5��˚{i���&�x��ڣ@�	c������ x5�0��(ñ<\m4�EZ��t!Y��k����3�Ro�p=�8�ө����uK����r��*n}���|Xv��8�`Ԁ�Q�|�C��Ȁ�f���_�SO7�/��֗�Հ�a���ZF0��r/5_7��]KM�GP�Y����H��Π�ġ��1x�����x �[1��KL'ʘ����X��y�Zry�a3�ܹ�?pK>�S�eι����^�cN����vJ���{P���&�'/�J���#�z1;������V�������TMݼ
5S�h>����V�rQk�~f	^*0�>Q[&y&���?���S ���քQ/{���!����(�X�Z,��Ն*������q��5r3��B蒨9�c��cG7�T�/��>��%��?����5F�!�nio��o��l]�w�~C��s�{ezg���|F�N\:R��(�M�[ͅ/S�s�>f+�y�Ж/�D:���v����Tb�~1̩a�|����`'���bz�
�#o��ё �`��ΫZ����}��L�{=8�������(E�W�_.^��n���uK�hm�� MӶ���>1��-�Ȭ^�ID�O�,��=�S�|T6ђ[��b�_�	�!� 7�_���]E�N��ȭ���Ym�*�|k�����˔.W��;U���J���t�ꀂ��:҇F�5߹)�1VGx���nݢ�R��NAkN$���c�p�0�����ƛ.�
�+��N�D��UAV)��{|�g+yq1�+t�pKZ#D�t5�ͼ,��G�E#v�}�9��!�{�����xbX�A�\{lJ�;G���9Lq~W7�m��]ѹ%ø^�����	[Wv�.����L��F��d|i?�k��*Rx��l����{C�+�ӛ�a**�*`���$�R�k��`��`]b�ϐ�,S|K�*L}I`#�����g8�4k���tq�#�9-�W	�k\��]�8�RJ9��A'�B��z�;��0���M��
rZW�k~��Mp��C2���ߋ��qR>f$�;�{��.��)�]09+|�U���6`����)�&���9W����1�5����T���ɺ�UK�X1v��0�֗F�`l��f�2(Ϩ$/�Ax0`ѭ%�3@*�yK�g#"�����|@dv?P�* '�����d|�j&0��=�T�zbR�N�����!*��;r.�����C�%�������Ad�VC��^kI��^��;{�7��j�^2y2S�D���lI`U󒪉R��¼�ӺؽZbQ��7���_����<z���~��籼����_�E��|�)�1G�ٍ���g3vw�3�0|�BR���VR#���Q4T��!�}���@����,���K>
��y60jbt.7�X���^��d`
���	½� L�<ᔲ�ۭ�����'�mr W��P�<���]��y��BU��6J�1' ("��_�z\���a���6hO[��([�t�#���s?���fR����l,߃�#f3��{V�j_!'6���ٸ�/���1Εh��]��G���d��5�����)��5Qi���by��٢+m��j-ГU�T��g��b�p�ے�=�_W7+����,�❧L�3_���=���4';_s.%��yRM*K���� ����\v��Fw�	h���?y�,�|$�z-���A�4����y�`�
�<��ph?<=A)���A0-���XH}��ip��>��xa��1��2LJ�#Q.-ty	�8�����%�ph�D��	�N,�	�NU� �ú��Y�V`ë�T{�O�y����>3������j��-cK1K����BN�8g����
V�H4X?;�~f*
i&«YTlt�N�S�w�����3(O���a0��v�������w�+�ޘԫg��?ϝF&�h	Fs��r �A�wyǌ��ц��)����؜�ۑ�=O,�����f38t{���V��SmI��^$�+<�A�3g����ȔYm�u�6N��q��yh����y����GF?e��s Q�xg
Iز���d�7_�%��bk�4�_m�[H�|�܄{�M�R����՘��ك?�w��R�*�W�#�
�I1(q@�s2�6?|��*�R��"�MP�T�>؅�_�x`��}��\��	��ղ����-��A�>8b ��u���G���о���
�]���f�����	�͒���7���V�!z�,��`؉0W&*���]��	��t�  �㗄,�7 *,�5��ko�8��� k���bc���il�*��gt;���*(T�M?���3�]J����B�1��\z؍� B��=�� ��N�[oF�$��t��f��N�zSc�>�j\��Z�qݯRY����J���Q;護$���>�c��g�et�F|�s�U19��7`���P���|Gh��� ���T�B��]}�7W����X5i2S�n���騭�&�4����|��"���(OG�7IO�s~�;��Ͳ3���(O;��}1zGw����c*.L��.���`�=���Ռw����H"k�v*״{�o�{�Lnt44���;Ϻ*��)E��`j��Po��2/I0��O{E�X���!��H�>��C������K�Td��(1/Ϯ,��)��A08^��{�+-�.~�d("cЎ��N�5:��)t^E$&o�}�����b�����D+�,�n�$�_��8�qqt��>�����e�=r��t]�KV����=�����R@t&�l�h+H�"�-�1&���.�����E�6��-�]��$aͣA+�)��Z��"�}O�~?��N��Y�N�d����f���1]��������ӻ�[�Q��څϨFiy1 sOjA����Q+�e-b�U��ӝM$h�N����u�*��|������n
~l�QMqg�(�
�y�>m�C��`ץ|I��r^å��f%�����V�p�(R�{Y�vfk-aA;�c��ə����'�PFJ�~?1#�م��s���m�܅{��ZuD*���H����e�:�tR)�����������
x����&[,K���~�Hf���n��v�"��čH��S#ī j/d��G��^�t�~t �;�O>����@�I
2�I�`K5�p.���M�VA����ʰ�r���U�l���-��;B��2&��=���l��D�A^�V,S��%�F�\��4�}c�8O���O*�E�If�Tds�.��TE/U��gW+�C�Rc���� ���oEKS��Cl�1��iid'�N=x���(�@;�nu�B�6�N��..�K�[�� *'��h��7/��u�9��V����|�w�}��۫��*)6>��D\P+��%�&)z%&�x~�,��-Z�Ԍh0�9zb�e���/jU�,[N'���6c�+F�n���YOW�pe~o��� RT�(��Z�@��!�#��&�pn�+�z�P��I�i|\�
��"���U���,YU�R�n��fP:�D� +����*�i%ͬT&�mo:��P��:Z���2�-!Ƞ�c i��m���s|�N\F7�e�@�:'���34����H�ݘT{�Ӫ��L��|P�cff�HV���٩OWN����׵�U�E�����1I ��xa���
觠��t�R�h����=� v�ܬ��O:pyh��n:�ź�m�.�� 4i��3��� �������u �Pd'�נ&���\V.K8��
��k��A}n&ΰ�Oys�0�� �� yꄶ-�uh:|�8�`��\v����B���k��(Nt��F���B�a]9�ccM<ȿ8��_;z7�$��a�.�98l>�pT��[��x��!T8E�YJ�J�ݪ?��ڭ���|�ߕ����h�Dؗ�դF`�ÁJ�d�G�^Wʙ�8kb�M ���n�Q��x� !C��D%�ARaU��8�h�"Q"\+�Ns8�t������&��P���W��rR��(�����c�;�i /�Wp����k!��3A�j�)Z" ������CTБ��>��h^g����Z��Z'=\?&��!L��
�~�Xy�� �,�h��1����YI�|5�gdcF7ǭiG��k�Y�n'��{C�v_m��qRu��}F,+�[����?*t��gG��9s���L����	����J�������WYd�Ѥ&��P��q\�~M�T��ǩB5�{y]�B���A�N؝ޅ�Y��W�(GVd�q �c�u\eP� �5�_)| ��8 ��6��Eb�Z�v�ٯ��Y�+���0 \m�s���d�ǘ��|iv����J�y۩{n��*���+�~C̥2S����Vp�Ia�ߣ��z��kw�gkN���L7k�DDH�Z0!��Z���ֆ�G����Zp�5�oZu�;���?��m�[�gᄳ���[����+�R`ڙȔ�P?��s�F�I��f�3��X&�Ө�+Lw y�Y+`��9�;<ŝ������� 8�	-b��r�6E���ܪD�Ȕ��|#�&�ҴS[�p���WHJt��_'�s�Xӯ���KrIf����M���mQ���	��}k�]��ZJ ��u8��l���2�=XTn P��eJ=��pT�؈R:�-�N��~�7$%'r/,l�>�@�9��;26�t�w�{�_"�	f�f��<����D�dM-;��ey"GL$z*�)d�u�/�&�
��p��9� �!�0��"�gc�4���nݡ����r��Tq׆Vl�In�)��tO�b(=O����)<h7WD#���xdM�R����+�'����"5���)�4r�R`��}?�v��n���D�<�^�2��7+���HXgֲ�%�F��u�Cr��?��}���~?�J�Ң���Hu��=�7�����9��1TՇR�دH�PϷ�	_u�~A���ֻP���i���re�IM�o�$4�YAc�--e�]]��/y��+��%'+��u\űyI�I2�3��� �߂���/��>�ъ.�oҤ��/�I�ܴ�OF�.-erLǤ��|$S�@i�)���C��j����DI���u�����><H,ْ4n�0"*-�"�ЭbY��٫��c{�f�7��[Ѓ�ƅm�Watɍ��伊lzT�D���89�8�m�=��T��j{���Nbv�6�:ZM�_���}�{�,r��	*ǔs����%a��o?_7 ��$z)L'�y[��ռ�0�'����N��Ң̥;<|�3�EH�XB9@�_��8�b�L�e��m��b�'ʅ����G5Qڌ�_��nX��ap��ғ/�XVs(��}�3aZ�l�~�ʲ{���}�x_l�����R��wGw��\w4?�K��-�N��v�4�7�< nHT"�eI�܉�ԃ�����}�U�*!�Î�b'8�|����+%����G����U��d/)�lr�p����1jCO���(·�hJ[�1*L��T��Zh][7�>������+�cc�c����)� �Zҿ�Tu�����ɲ�����B�<�yD;A����0��HW���)�q-�Tˎ�?XL.!�~Z��_wʢc����BG���w��G��׵��y�{�x���"'pҷ�<�9����f�����@iX��4$�ԭ_Q:r!��e|7 �6�v�����5e�6]��Q�ݝ'�p��#�l��]q0��0�Ӄ��kX�{'GTphA��H��*B����Q�jPTnd��B�\��*��n� +�:s�QHQ�����ppVs���[��P�u�ul�֣�i�-��N�?�6��b��m���
AA0��4�t�"���2����c��y��)�¾gȽ�*�s?)���b=���}�x��'��I�lu)��_s�`�M�b�Tp�3������t��=��!�Rc�F���ڐ���bU`�^h��[�<���?��PR;���Y9k����r�n�^ǠPr9�j��d�ECҕ�a��|hnC1�/M�*�F2�⿓M��ts��0�o�D0�W3aW/F��������S�q��Bn(�w4��-�v	W#��K���x3��ik�L�������c=�2�O���ۙ�P������_ӒCh�����ܬ��*E�� v�RW?ݣp_�*��?�v�|Y�JVK��p�/;s�Eܙ��a#i��q3BB�.G(����SQ;4��>��6�9Z�uz˞������uI=��\p�B@l<,�H��az��aÜ�9:�2�Y�����"�coy�ء �����-����9I��Y�ζ˂
��T*��DF]�M�ז���u���B�o|��*>���"���[4�04!	��#5t <�I����_����Fy�^�`�����-a ��w,��t=�$�~��`�C��7��l���Uo��;x���w�N2F���Z_���Q�.(�<'d�a0��=P����=���>!�*��~V������Ճ^Ƣ�{ʿ=��<K��KY�E���K{`AZ2���{�� ���In0_U�K�����F$���T����΅9�p
3�����j�\#�g4��ty��L�=�>��q��=��<��l�_ˍg���m�4��GȾ��H;��#Nl`2dY�T�㠊Vk9��nZ�K��	�t�į������7o9ǿ�oY{/h[Kť�,1��"-nd|پ����U�tp�3D�/t=��q�����JD:b&(
.����eBǅg�np��	�D ,�"@#f�>m�S/i�Yt��A�~Z~����i�@3��ȋFel�b�*��*����s��z2�d����n��z�B�I/6���������A�.U�1?gG������A�0lN�k�)�lN�ĥ����:E�v��2�n��Km�8n��b� �8#,�
u�|�,ٖ,=}(2��΁%[R��zK�T��{XҔ��p4�
V|�^P�;�� w�Nr����D�����j`�ag� i���H��9�%Xa�r�r�
�A�����u��Z�L1�Ήj�D�O����+���X>1�Q�p�0�^p�w��z������7�p�H�:����[��5����=UH�Q��X/�_��C��Ք'���v=O+��NT�Sْ'�#�㹫�[ �
�SV�$��%�<9�zf����2.C��\Gvl�������>�[ɲ�s=����%}���8�+�`'�|�������r��8�4!��n�/�p�ne�|����&��ظ���(�O�M0}����/0}*I���d$~I��̨��n:=!'wm|��VN��^D���(FIC^?� [�4y���R(f��~?I�����_q��=�� �_��߲s2��
�A��~�,�6�+�S
ĸK�ė�����tr�ᏋR<|��qno�����e�a�;�=���7
Y�>qҀ��L/cE�fr̛��q<����4L���Lnڥ$?��<5�ӽ;6�BQ� �m�dt���ġU�v� �U����g��m�a!B%%&��δvHY�JKMw]|�����$�T�Tx}�h�AǨ﨤��-������[w���wZ�]8RFn��3��7�o; �LT#����������K���(�{�Q~`]���qt�|���pO�\��p�#�%�{&����\��hG�Kڗ'=YɠE����I�ź��#�m!i�O�3^��Pz�i����Z�U�'V�����ܰҏi�)���3��?�b�p$c����2��&�~Db%�T��围5�(��`
���M5� h�ㅶ����P?�Ɖ�&��5��Ξ�L�S�y��:M��\�.��Z$F�Ͷ�4�f�Y����'_�H��R�?Z,ő �gϭ�_Z�R�%k��!^[ӗ^�aM�ʠ�O��ekc�b�D�qݍT����J����qPOpi�����v���{�Lۦ���r|M/$�D�"�~EsO''��%l�8��\�27�<5Ҁ��lϯ\_���E8����|�S�8���Ϧ|#@�8��~&c	�]t�փ��!y��~ݣ��m8���`ι�:]�>�՚�/e�\I�I{܀W�G�@�v��;n�����EI�9A�fԎ,��ո�0����b�v|V����"n�$��Le0B3pvإQ�㖪\���5�E'�ua�s�_D�����/�ڙP��\
{�%�4s����z�p�h/���A�U_�Yn�.gY�Ɗ 0=n��.���Q�>����t���ޭD�-�N���(ZP�	�<Q�+&O�K,
� v��E$:�ű,TL�ںלQu`�I��%�G�� ���m�j,�	���V�rW��*$���8��J#�RL@�f�. �ɼ_BM�
3*Vr!���E�t@�nm��w����Љ��?�щSk$kGo�|V��'7`����J��-IZ�ɓ��3������@X ����g'�O�y^����'X[ �z|D�6�h5�G�U���j��k*w`�Ů,e� �F�<x(ƻ-�|��ǆ��������x�@@��/�5�*�I����s�7$��j���љ����(�7��W����>�*���ßDo$��^�����ݢ���-��P��T�e�����@�4���1q�y���\]f$s}	/&�&2��Gm@����4lOK��[I�I9y�]�vGXc-f�5������&ΰ���I����PH<�����K"z
Ŧ�P9���v*�'�H�gVl�.c`e-��LE#8��0�%�}���ʑ�s�n���~X���Lĵ1��J�cx�g�`���4�0���yg��U�i��o��������m{ژi"�K���,��5�a��ó�ծ޼�	1?My��n�?�6}�(��hyn�@��bj'ۿ��ZR�c��ϒ�qR������T���OV`#��&���c�aJ;y)'���m&F�(�l��3^$^t�;\}��/V�l�'o�W#d���� j��#�tn�Z����!���d���msT���T|�Ϳ����(0�{O����6E�6p�b�g�DKnN����s	oA��n�EBz�U�y^Uexf�a~��q�x�*퓮#�fnP�u7A���NwSp-M��'�g��T��;�D�c6��q��[�(�K�iB:C9ɍЊ��>��i�5�����F'�"��i}H�\ܛN0��� ���θ}�oe�2��s|�a��oM��j;:�3�JP�07�	��Ωgӷ����J�8�jmܔ�҇N���IS���ݲ����H���B�{�53/�b��M?���5t�"F��6���0�w&�\$C�� UR����D�:��.~�	V����JC�7��$�x2S�Nx�>�kV�_�A��R�<�X���D�O��F`�~~u�(��ȝ��ZL. �����t�=��"~d��3����߿���\1���(u"��cĦ��+��s�ݘi| �SAs��,0)����9�5�O}�f��c������]���A���ҙCI��4��J�߼UM�x��ρsDe��/]���Fw.��c�F��66�D���(� ����3��i���9���f$���O91Z;K2;^�]�+ǵ��d���	噞�p+�����S��)O��X���!�^�b@80����}��C(O|��R�>p��`D"�k^�ZE&r� ���֢�� Ъ�*c^J�n]�<���G١%&E��*x����=�E�R~�����Z2l�̗�~!�p��A�������/�t�Jpj�L�QTt�<�(��-�e�C4v1w{��Kr1/#���b������tʙ��7�PK��V��T�_:sOC����m��U�짾)˾��cC��"�����G��͘g^O�=d�.��F{X�>�=������ Z%@�C�A�nڄ�c�yb`�H 03J����QC�k�n�&�C��%�F��^�����Ը�Q7ͪ(�(]�d)їl�αlv�h�L�0��,+wI�!����x����@���/m� ck/�^�CZ���;�_�\¥�6n�]��1r�ĜO�������!ݟY�K�*'9��/Z{�Ƕ���8�g�@!}��4�\`�R8���嗘De��mp���F��!��F�B�,�!Ebs
~��WB��O����m%�������ω;�5�;�xE�2]�㟿{�1g;����u��N�({[���&mٻ���2xI,ܻy�Ly����\���rЋ���%�:Y]A�"��]ɜ��X�!��ށi�S�S������������nZ��RK�KgW�׾���Կ5gp������7�� ������a����g�iAO��5ρM��mӈ�8n���|��J6�ɵ~_�ĔLp�%>;�lg��,v�g�$װ�pq���G�����$��H��?��7����1Csnm�כJ����''�G|��m'��$�<� =E�;*�u\d\:�5�J��cZP8O���>y& B�C�|)4A��i)lN0%�lge2�ܫ\��՞&
ȫX4i����	�Ѯ,�4E����6����L��z�2@�����a���T�B����H#Yj�r!��ӈ��H��|�����830�;�==FZќ�6��~Ek�au�<�+<U�oK۵�A�5�d�q�I}kU�'�C�����<�� !��-/����F����ɮ�QYvj��nE��q���%�G���ᔊ��9|({^Q�J(7�% ξ�	;L�o�p�q���T�e����YX�l��3��@������`�+s�﹙y$�O�����:_&-9���|�Ri9��>�9��c:l��w�A�66�=v뇋��`�w��c}��E;�2�,��J.)>N�FT�Q� ;F0�2�sq�n�Oԋ
L9/oP�Ѻ�T+����v2ҫ��/�1�Ezm�FLyH�T��)2��=� v�1S�o��:���n��8P�P�~zQ$	),r��yf�A���eGn��#;�P!y��µѰQH��ue�W�W�Oܰd����`�,�7i���c����&\/�L	2����.��]P��f�"}r�z�U(��g���|�JK$c.�!i�����=Z�nphH���[� �/�����Hw��эz�u{X�:�J�Ҭإ��ϋK�27x��/� ��69���(Ԗ�����f�8�$�<��ur��WcdA��E�F��@����������$B�/������j�Qb/�eY�ݤ��6H=wo�GyYn�.��>S��<�l���{��1�A���C��j&f�;��E3�c'd��j@2���F�g�E���0���P&э�a��9��+�Gg, .�6:�{�[ıa8��X��&{�U��=���\[��Xg���
�ݪ�^G����̈́n�e}|�)��h�F!o�p�?P|h#�O��֭��{ F�؆��χ�47Geŧ�g[$�B�s{c�y�����H���T����tJh�5>�j��$D#X��4F��\�ydL�����3���6��?wy����l�ɤ�p	�Z5�Z*l-��!(��Z@����.:�a���`ܸԕi8�O��G����i ^=�J����5 &���z����9�[���5!��{%���-Bq�-�plVcN&�/ߊtt�mן��tt���V�+��-����"�d��oW;� f���2���բ��n�\P(Z[=����.�N��M���ֽ2���3F<vBUY��s]����OT�Sw���rLy�W���N��a{Z���C�_<~%/KS,���Ea�)yZ��|P�bltt��Y�^�r�H��O��;�Bd�d)�3���.�`C\_'XIW=��I��yY1��h�w=���s�+��fjN�Jtm���wy�P���a���x�A|X�	�ŝW|�M$�zQ��p7�5 .�{�+���X��\(ZK}gi����f��h�h��������u��Ŋ��Vc���Ex6/yU�wŀ	�ty�Q�Y襗�fd�u:?�b ��98|�*{6�L%��T�*��A������3ڮ;���T�M�}]�[��W��(��q����^�gxn_	
j��Ǟ�վ��Ki�Si�p��'��}��S�e���?+qv�FX�����3���`���bODʞi�M�������	�&v9�eM�(�.��VF���E���b4���* ��&�p"���ɂщ��O]�[� ʕ>���j;$��V7`��T�6�����K�Tt�w3p���P ����ރA��H���r?�c��OKِ�	_º���[���#\�/5@v���$��ܠ�&�O�w�������Uʏ^���)g�,u%i�l�( *��q$|w$��M�;Q2����E�NWd�M��~�c��6$�T�]�[3��}j�;��6O�K5��:m��0�/�����ց�{?�;���&�H�X�ȖH{8e��>��*������F��c#= �і/mق�����yQg�P+R��r�y�����$�S�5�~Qx�4,w���� -e�W��g�>�`I()�0�,|+����v�h�EJd��&�j(k��qI�=��n�.�����i� �˗{�����9��ODG��L�/yA2��u���Cf6P�Y���P�l*���2�G1?+�}�� ���⯕��@�u֞�U67q�e {��am�������~�E�Y0����9�0D'd��=�|�*�,�҉$?�_�C,����&i� �͢P�I���8KĞ/2���f��3j��d��o�p�_s,��Զv`ŽGP�>.L_1�	D�)Y��I8����_h|�|6hC�<[Q�k��Kϋ���T�M�y�"�P���l�r������1�],��'�K�-=��e|i�]��5KsI{���?u~j�ѹ� ��kx>6S�g��̂Y��i�<Pb���2��{uH�-���Ș�>V�	�6D�1����w}�+jH��:~iK.:_�̤���T��}�N��Ĉ���z����i �l�=�6�Y�;�q�+�̸�nB�mt�,7�����U����F7����i�|�'��Dh�����Od���0!W�l\�>0���K%�a3pj�	��QP��%̴���՜Gk����`�xr��7�<��%�L MI7i�u�M�p�H,Ѽ��<nJ�N1�2��:��egaz���;ai�	^��9q3I'�Y�eȷ��:�s?��3n�^H��>���Q恡f!��p��:�M�O_��v��b3m���!�B(R���o~.��g�Й&o�1&F��AV�y�ً��qل�1�g��xT�{�Nl�@�wV�����J@Slh�2�,75'W�I�ʱx�uYbd,�0ST�2:w�a-��_s�Y,Y��Ý�F�����G���m�m<�uI{��H]��:%�$���zV��m B��2�&G�C>���h�m�����9����|ˠ���F߸CޚH��*�<����Jm�EK�XY���3H�U�_k����=z"!;" ��L�N.�9�,mEⱯM"��ߌ���S���F}�AJ�c�&Ed�����w�~of�*��D!��P���<���؊��&hD,�ɬ}·e���
4�p�e0a������~؋� Sql�?�`����tޭF=���>�c$"j��*ue�-��:��C��Z`��'�N�	����5�8?ix)G�.�ğ%~�Ϗ�O��:l�W��g(-��i�)=��;_���������;����S�Q���H�_�9��w�Z/��|Q]�A��#(A �4����WOy���B�Vg?cP�He#���G���)OZ�^ ��.}3�ݭ=R�?J�g�9%l�7�Q�� ����[-��H��dۿcc�|&�E;M�|k,,�ؽ�m�ȷ�� �K�M�l�Ms>��R������ƩY�����<_����Υ�M]fnجz��㍖{����y7>~���O����֩�w{���|�#(��y`�=�.��
�h�Q\�P��w�����P�G��E��1<.�w�D6vX�I45�i;q�m\�(9�EO�6lbAP��,A�>��U��us�L�EU�D�=�m�u̜��[=���K�6W��5/6��q��Q��^��&{��p���zҵ�CEW3l2�9��}��$?�W�e{�d�0&��!-�&O���<+��w1�d�L�'֌���]'.wq�fo:�+��1��̀7����1�\�LG��U��w��{�اL� �7�����?�>@�hy���&��@znW�2f?aiX#���������v��R�O=�X5ϋh�G���Ke�qu�^��^�aG]����$%f�g��rVڽOk+艉���hv,5�:s��`�^f���-��1����P(�.���}ե�i����][�Օ]�aC�eB����*wJ�f�S��Fx��e1�H����B�\ q4z�J��'�[_��Y'��hbW�o7��6�12'X�=�!�l�j��lX<���}`.Tɭ����Ay��i)\�RvNR���<�1��m"���!,��OBjk���{("�HH�� /�������$�P�p��.6�G���ף��i�^o	��~mwZ�v��=�
o)��o�Ha�@�?�8�k��p�S|-��G�bYҡ��O;z����/hP΁��O,At	�����$8A�[1��"@��J�e�L5��Qx(��,�uEN�٢p7.12]��w���W�;����NN�KyCp��P3c�=k���Sl!�z��xs�E���ND��I��v�Q�^�r�j�a�+�j8�m���ӗ��R����LNZ
�������sЫW�Q��1/��nBT��vO��UDxQ:)40�vlbE�I�
o�g�'�ۧ?'t	(2ȴ�]m~�'�7p�嗔���B4�{��T�����h����7���FsD�B�i�\�1��]������#�A�G�5��k�k�s~*����O���7Ms����|��<�=p�f�F*�~?�~b@��6�rLƖ^�#������U�^�Bj��,<�Q��W&7�]�����$���˭E�����?�{1�6⡪��@��e�^�͝����o)l�iv'�t�����;^]�IA�1_��[�(O�|�D�=�iɎ�#[h�`����A�J,�7bW�|�d��?GK�ctF�&L{�T��h�`�2�����_��e0�a��t�<Ǉ��c@��@e����y�e��°t��1UP3Huvք@���?u����>�W@m�<*j>��J���9�D��b������޹'�c>�2�D��G]���+#��5�R7;kO@+��*s���*qO�ڤ*������$��+���:!u�`x�����>��Q�'�d�R���� ��㝴/�bPS��"��ɋ�P
	�zh�5��r����2o�?RC��iY�G�R(�+��L��yRq��3�@���P�c|	�9�fY2\�Z��.��O=9�F�� ϖ8��n�%,�} ��u��^�p�.٫q�>ee��i*�I�?�����,h�����f(���d�������.'n��6�:�^Ϯ��&�����_�v�P)M=�U��#�FS>���θ�3+����DZ8�ڜ�͝�<+ܺ�g�Wv��"�%݌	~h�m�G����������?T'� �����f^Q;�P���z���:~Dwd�HK$�M!�<6H��^JIі9��|w���SW�RT���m�!�_lᘶQ�䞸R�෱[%��(��%�p:��N��x�u����S��R^%�_$�~����:5�2�QQ�2���(�v|�OS�v�4�� Q�P�rv�W�G��攽��"��Y��|���)	��f9�o��s�M��y�F�����dg� ��:����|V�4�M��Oþ�W�~@�g�>���c��Vyaf'<G�b_NZ| �j��k�ԝ'�g�)T�OǞ�t�?���B��2�t�7����xA�+��v���ZXv�e�B����z�#4�x�Q��&����1����:7[r��K鏲ẁi# �j�y꾺?+����|�;��:�7���y�X��d��F�;W�%�
���^D��R��{S�� ���ZQΧNh�r��6�s��d����9�:�<4�c����Y��(%�m<؆ܘ��GҮCK�4#Z�rgFU�˲)/�r||(�K"�B�����ҾH>�,på}���o�=n����W�-9;�{1�]�"�i\�q��t���h9�`t,���O�+��Y��Oa�{��,���'����<&��ֱ�d��Qk3�x��N4�R��>�����c���R��M� �@���|�8Q7����jt&�����b�(z'��h�����f[Spd3Վn���5�G��/��%�x/W"O�E>��N�T�?1PXt_��%01|X��L�b�=B�s�[~E����nË��nmG		�o.�KyG��Q��q�Uq�QaO8�6ĭ�ȩ1���%��W~E7K~n��ɀ�L^'��z.�:je|p�S�F�)�BP�c���.X�J��?�L���U2� � ����^�m�ö��v���:/L�:����_��`E�F2�kV�a��*����Y���������Kg�ͭ�ohm�פ%���c���?t�����3�5���2�`����F��2e*���^=ē�q�Xȅ�:,�� Hͮ��%�0E[w�b�-�6�{�q�x�i��]�a,�!�p+K�9�b{��Zx���\��ۄӔk@��m#j���)�$Q1&�̓��l���<�+5�lU��[T��V{i=���,����4*O�Sݯ��}�a*�NB���P+��%(K�V(����<H'�p ����<������1�l�>HF����Գ
2Uu�pNY(��M�*�4�&j�R�#�h۵3�����V.\�av�?�B�ac��<� ���{*M����-�p\&"��d�#���g�L��P[g-���@�k���H�0�Oʄ�WFk��{��	��/�%���%��T���S���R���'�BJ�X��hR.-�"�����$4��P�<m|H�m�y�-��Y�>+gg��o��y�tO:ڒiL�t-��{��o�s����� �ݏy,T��-���XV��(��1�R�?��V1���ڀ�9�\רt�؄��L�Y��6��/&�d��#���i�GBȾ5Y;�$���������ئr@v�x�Y'�S=��������u��!����wւ�]+A�7|.��i*�Ox/���n)Ӡ�_��K�a�f�ܗ8�{��6n�Dz,%h�P��D�䚘�{�"��V�_à����t���`=���b�'�[��;���ݮ�T���^mz�)�Mn0:⡎qy�,]���s�aT��6ځl���Q2�������3������o�&�55I���NQ�@�3����M�~ �Gr��WD9M��b�^`dn@=^�C�����|*}���OsӈWZ��>.�bA��*D/}o�*N��*4X��ф�*��^6����<leR�;.�ʸ�]���:+�ѢB,�&#���]��3*��L�}8��[��^=͔Tvw�y�;j����^��i��������	��3�4��w�mq��oX�ʬ�,���7ſW5o����{���������7�+k����b������8ć�'�6�ä�1���M����mkec&1&/ߞ*�e�X�t5���3���$���*RV9G?�HqS����ڌq.�xyV֫�c�8�!��	˯%%�r�<�5�\;NŴ��������w%���J��T�X@|�|7�p=x5��ߠ���m�?>�e�5-B4 bQt$��i$��6�0���6�ز�|Ǳ�:A�=y��!�1�P�=Z:�}Ƒ=6kR��0������ږkmd�v�����O�; �	n����i����3�j==��_>;��RJwuy����f�g�tV*�|cS���:[�/���M{�����ߨ�� � �'���C$
�&qM���c�~}	�ahDX�Ó~rf�Pk�|E R�"aՄ�\~O�i0k�/E�����k�늰��5?�D]�S=+�3��Xނ�sr��B�F��-n[@�p$��y��o���6�����L�J�D�lڢ�T���iV�g2u��6bP��Py�$f(z�;�k�����Dq�}#�o?���W�l-�6�-S%lR �(���sL��C3n$��N8�\�s����slc��a/�f�n^(�r;]�\{n�zE�k�u�7-���UX�&3q���ih�Z�|:�\�g�+�gg���ǟ�>-�t���q��|zBK`��X�t].��r=t�!ҵ4���~�ڔ�4m�r����\�V�ﭻNߣW�M���de�pJ�,#��9� �L�e	�i3���]��2�ĭ�l]o�m*�7 �d�,�kd�	�xWX�z`���Wl�b�L��2��]�S�Oۚ�N��$c��w�|���wA���X���u����5� 9V�1o��F�E(D�#��2'����	<��CN�?�NF�� &4�N��6���`�������SȦ��n��q��]�֖ ��ܜ���ی_-�2Q,:+����ɕ}�ݭ���2���g�6��1����T'�}�����O2t��턹vxƈ-\H�~�US{���=��ܮ�����P�����w:,��VQ$f_��L�h�nD�@t�7B/q`h���XE۽kťf��!W2ך�򄿈dY�w_��G,9��AW{G�#���E�,,+��W�g��d��ΰWT���)�h#��ro�${�?��8N�hO����Ƃ��OU���!����PfuL�~Xuk�;Ȍ:a���16��eLBfg�`�$Z�����DO���[F�rE�l����W��1�m��9�h6r�ۘ��%!o���.#�6��=�6[���tt����~~#d����궟E��t6.�C�@.�bv�m�\lHc��2��-�~j:kNۖ�bd�uM��{�`�p�j���	@iJ}�׳Gb^-_o�oi��;ޭ_��2���b�;,q�D�M��^Ic��}Ov\dipO����<����ʅ%&/Ek�%ZA�"������U"�~���1(�䥩p�����t@�0��Vʠ�n�G�3	:�G�Br�og�Þ�x�k����SoI�t�q��7��G��}jx��u�8�7�GBk��0�>C�{�_��N�O��Wh7�[v~$�b6��zw����eh~?aQ�{�t�\�?T�ph��ۢ�QsډjPd����b}�fdl����S����ū�4�&v8���B��ۋ�J����۞�=�F�b��܇�����u��89�a�6�ny���q Z�}�x�N�L�r���om�>�I�,d���P�Y��:sv���T5��%w^�Pۑ(�hg�4��h��X����<��,�	��?�+�P��	6����\L[XQ��>�G?_M�\��LtN �ʣ
�|/ö-#��qV#��N�v��7r�;�ifIu��v���̽C����}XȖ&@y`I-�N���]]qpzlw]��g�w?1D���r��l���	�E�Cs (� _
8�<�Н�0SښW=A$<��n���$�i;-o��䭇���P�L���*�"�E�[-�J����\��Uc�ge�K FI���m�vzh�r+���k��dc��N��K`������_3��<qPʏ�ݏ��G����Q�u��
��w���c�G�F�.��)��W�먂��rYj�<�$|[�����UO�&����� W�D�/�[�_�:S�r���	qG�7�X��/�Sh]Bup%ĸ׋��Eʆ�%xd;��kً��Vlش�2����ҝ�m��k��rzp;���r��㆔�ˉ�{(b�Q��mq1z��Uy�t���#����˃]�.�ܺ~����ӲV����h'����GD�7�k��S����w�����Z�U#������(����#6]�q��
yRm|.�m��ŕȼ�稆?���s���ᑮМ ��d,*��*����F�v���A� g����G��Vډ�&�6��ҕzn�&�r!��h?�t3	;��,O�њ/,�#(D3���4�l�Mx�,�n��:~��4��r�
YkP�+�=*�2v*���`5&������ J�K��|K@�>V�h�< ���sA��R֒�(lW{�ѳG�6wFM��%~��8���K� �3P�)	���G��<~���� D���v���6^>�t.���O�6�Cz��ߓ~/�}�@$j�t6P	�f=�]��\ xDZ��+ۉظ�i�|���	w휷�@ۧ~�db�z��N���2G��5$|s�[�*덋��rL+��ȅ|3���#�Z��u�Q0�dfǆ7U��D���a��4�H!4��y���P?y�'�׈�UH�H���S����2~0�N�q��RB-��p3�z
 hC��Ak`�TꜾ�Qnll��ڠp��i�5�y6��}]+�2j�d��tfR3т��bE�)S���|��#pEoѸ���CX��zx��ь���M��5�F���� 8Yk[�����h�b�$E�wP�/�$p�C�n>�k�Ǌ/.�t�h'����*�Mf��r&�*d�E��B�~(��KBCh��P�J���M��a� ��6�6�h�~8�p�i+QUqTߐ:��e�M�ZE�S5�g�.��^�m

�zJ�����Jhs����C�O,5����'���+c��k��~��
Ƞ�Yv�W�y���;�Y�`a綱��ٓ��2zg��8�g@P��"Tm8��:gU���}��$��и�×݃���NO�H�Ѝ4��[��캸w�U��+P����\��W��ɷ���U�NZD��v��H�s��2�J�A�e~�@��q}&`UUaY�5Q�E+�g'Ԗӷ?qH�:��_�\��(s��iI�۲I���*�*ѷ��6���,"��蠫��@��[Lfw�i�F�yf�����ǰ<7����@>�,�uf���kQ�������RW��h���o�ʨ:N�jP�S�c!B�����3A*Tx�3�4�Y-sM����ف).����?MN_� A!���"B񇷮��?�����!c�����튆FQ�1��k0���f��= �xR3�>�}Y�b/��N��?��D�vZ��r1pr}��i�.�VK��Z�*�c`:�������܁s�xR�>���*�)`��sK)A���战E���)^ p��+�A�H_�L��-Rp[�G��H:�=ۈ3'��җ_:�ah�J���T®�[��)H����{ҡ#s�R8��qH����ߋ�5�DED����U!��0a�ʪc�C�|z��|A��D�D��_~�������ŏ���Ws��u�.;x���/4�RD�Ĵ��0��q����0����Fk������#IN/�
�;n������j� �W������M�5C9&\�'�g������Rq��'�l�eGkJ�rL�=@�R	�ϊ����Gú�K��p���5ܮ�N:"�Km������Y�R6���~/�p�����mSE��))[�o�����ׄ��U8�����0�I��N���yNV4���K����춳�!��j�҆a�:4�N5+\���Ƶ���O��,��hv@-�`E��D�5���)g�ۭr�
&��niً
� ¾h���H���"R=�*���r�R��ic����]VȼV.�;2c-������As�ۜ�7c�X�� �D�f�S�Z<����4�9J��w_[�R�������*�vR�8PG�uxi�29����#N*�`z�j���}���m�邝�1Y�?�������D.�F 5�8U�}x�޷��UM�Q�[���~���٨GCsA����gnm�-	�Ű5�������/�
�i�ݣGیn�l Q��Ȉj-wʔ��8�j0��9q�1�{*-ρ��� $��GH���
]���-�Q�r�d%k�c�zٕQ�4�8d�A�Hu��G�{}����	��^���f��fL5e"/O�S���� &�1��:c �|�ֿ���B&�M:�T��Uš	��cA�W�}}�Q*N��n��b@��҅�CG1�����v]�8�4I��ht�0)v�CZ��Y��d�h��� O:��52,x2�~�j4C_�F��@�a��YA-tȑ��\��h���v�ё��`�Ma_���.�����/۷�R�� �1Jrd����ܤ��R;ܫ�֑:�n�`:�.��N�)SH�yR�aZ�>�=��u�M֊�z��t���g�T�ݒ�J��A��n��ì�|m�T���W��uv�n��<2ff��y�	��k��`C�)����C+�����L��$fe��\_��f�<�m�`�6=\�0e&�"u�P�ۭ,�\r���~J�ێR��;��fɵԨhF
o�̾삵�!��U�}��4��eF�Еyio%���&�,����t!�"��Q���L=�z�] ��K�Q�h?��
VJ�SY6X��gA��0<�����Q�v��ۙ��\aD'�	��O�W��N8D%BϜХ� �4"p��r��8��߿�	JN�H]���`����j�7�i�7�.O��2~�C���_냝�0?�'@ҹT�}{, ;l�`��!�j���!@Ɓ��[�.���_;𘸐�yHrwj�!W�� X"n���n+r��L�z%D$��g͏��D8�����=T\!9��/_ [�Ã�F��'�oM=�XӼ��\/�U��������8�s�{����}�*4�\�ګ�6S���Vw:M0 ����8��c���
�*�&I�@;i� �բx5JF��+�E��PE�4��~3dB:Ͱ-�GU����K��պ���wct�).��O4 V1�&��U�{�ꀸ:ɥ��޿Hu�ai��N8���!5��D�U�7����^�E�釠w�J6�s��;"y�4����f���Y���C�#��+KY=�S7ˇB֓�N�Z/�h�����)u͂���D&Wz����X-��J}�5�<tݔ�8l`�J*kTx�<o�E�<aq����V�����|ƺ�׿�:W�7f���U�?��2��i���q��x'>�� Iu3
���o�JGc��ZlpE]5I�>���$���4i+֞�v��I�2�G0h�n-�S�յ��hI6��\ߚ�c� ��~�6��>��:h]qo����}�iM=i3��ʃ���`*a�
V�0W8ٲ,B76�Dx"�	[n���~e�ƌ
>���RyL�Q��pO5ϓ�}Ų��=�`�!U�`�t��+e��ȮΕ�ge	Y�!�qJ7�_r�:O��4a����
Q��i~��B��k�而�̔S�R���Q4��c����hP�z�Ǥm��3	�ۮ�h��&�d3�eC%��ζX����\�GR[��l5�9|ϊ��06(�d#��
�X�#f���ƀ�[(mHU1�����9˓�������+BR>�
�+�G�ն(�$�$�W�ќh,K���q�3��Ji��q8Y$a@b��H����n£y���J�OqU�bdMK�,�Yf�`���Y߫�����x����N�6"�v����a8���K��J{_>�����@P���$��5�GO�ۮ.Q��=�\�c�������l(�2����IQ���	1Hw.;L�<0Y���%��ή�Q��Iy�O�[�O`v`2A����CV����O4E+E���r��F�A��v�H�^��0�������T^*�{�CM,g��p�P��!��zS�Y)\����Η�d!�➻\b�����|��v��v��i0\i� ]�=�pC�U��uj�B幛�d�mƵ��f�Z0� �H��g@�BA!p�M����"�m�L�o�	�iBb $��W.��C��o��D�c{�,z�K[X�B[��?�_���rWW�����tF�Z@��r�Lv��i��t���(e'��{�o�e̓��h��!���M�����W�l<�u[�HtH�;UK�.�T΅�D�d�+-ϚX�xJ�� �sͥ�-�M�{�����*��qt_cglq�,qO�7$��BS"~�`E���z�Q+����>�Aj>m�e�GWG�Ңn�/�Z�?�����ŗSj�e���ݣU�Mխ?;�=��a�G���J�����ܻ~�9�������B�y�O��#�*�m�S�׿�D!����wȹ�8��]�r��1̖���ך�Q@9�쿡��D]:m���R�9u@=��T���rb�Y7�-�<:sp)����+u?>�_BI�W�Ѫ��>:Giz0��`��SQH����a�"�<�B�a�ӊt�`�ڝJP��E�c�n����9�\~9�k�ۧ'�գ�B_\^8hL��X���h������[1�1H�h��������W��	���@R��0)F#�D(I:>�K��pU�B�gR�W+pBC�
Y܆�&/��rxn!�Ҝ����4.RQ����*SZ�4a���$���A�%q"H��1q:+dfR4Q�3����~J>nG@��]��ةG׫_��:�܊7!������4w�!^2�o����޹ѡe�q��(Ij�V��h���L���8ɟ�@��DxX}i�)��g�m������݊SO�r�V�P�:]����H��M�u$W%�N��RB�i��-�����U��}���$�GӖ�N�&��a8�6�b����N1�
O�O!�KȊY)pL��X2Dj�⎗ߪyE���!�+EMӈ����Z��g"���,8po�u��<�A�����8���K8%�G�[h��!�kg!T�&���z��p�*�8X��D*�t/m���S��s1-՗]ip�Ko��X;��;�)��l�Af�- 04�g�+^RxJp��@8)�HZ��,|~	ӭ��{���=�Rp2��|�9_���"������͒�d�ŪX旬%=��rT��>��[~Ԍ��7��Y!����x�Ex:�֑�e���N���Do.��]Ç�{��[l=����	T�����V!�����1��SQ��O͛�L���3�Q�s֠�2��o�e��(��`+)zȓ#�M���ࡥ��@�y�5��!����M�od6%����q(�P�@�����5�i�v�P���m˫ڠ���9g��J�Q�D����gLM>�G���u��</.PC�#>֦�~�Y�g��qi�3���%'�|K�%p����XP���	G*��L�#�9��a�l��d�Q;wٖ�r�#��e�j�(W\��e�R�O7b�ܠ�I�v������4%�n#B\k���]��x(���D�o\�,�i[����5���OZ�!�~҇g������{Isk�%8�B�����94���˨7���g�}�FNP��D��&,d�b�=��<��0�(o�H���f�?�>7�\b5=�\'Va�f{,I�	���1���_��7��e�_�z؎�9�2//+��_��/�Dk�����U8��D���EKK�d^Z�˷sI�|pAFA�+�>n_���0_n�M�8 �d���3���	�HaS�?�v���O�ީY0�d<��LQW�è�V��­�ꛠi����<{�6uny���/D�6�&9Oc��$O8�m,L�
�1y����I�����
�ȳH���C�t���6v41qYo>�$�Q[�R�xPOӗ�-ֹ��5ƒE�:��w.d�~��|7Gawh��^=�n;=�ID�_%)��#�2��&�_"��kVnL1�H��^n_5�N�Ew2�cj���8����\c�����\��w	��%{z��� <b�ƺ��	4�x�U��5XS�ni8����mܽ�}L��.=͋�f��ط�����r3����s�\�2��E����^m)Ue�`�~�g@�e�2�f'���~0u�VOM#~�LY�9�9�i������u�?�_������蝮}/���������pwU"@ihF���D�||m�-ͷ/H����3k�\����ж6������H�-�T�]59l [�$unj3�q��2�tA�,4�i�4���G��\�Y�* ��@W|�Y���^���R��Z]�rIx�Z@��^�|)�~��ztyA�S�����T�Z� �7ۇ�������KP�̸��O��#��
Xh*h��'�>Y%7�ݪ
9H-X��A'hh�=���1LB.��Q���J�m�U��]鶲(}�X�64��|�Ep��)7�� `I���=LR�����,�o�*d�v�K�AP�����l���A�@�N���x�Y*9['{��_���IY�E>t���	���ƀ�:�ʴ{o/���P=A��hz�_'���c��rS!W�B�B�ה͈%U�혷//F��@��������x�T����V�D��$J�� �/�S�y�[a�L��CgƮ6o.�^5z�F�U��\��)�8$�5b�6�,�])J��lix�0|�B�E�q2���b�Ⰵ^r�
�-郘���=�~��HޒB��߉�x6����v���3�L%x�����RZ�.؝8f�ĮAx�`y�#LOl�;{����w"���L���R�/��a�T4�Y��L�J��O�ٹg��GV�Y�!�[J;�Z�k<"8�X.Z���$W]5�t��e੊a`Υ��k�m4�n���ك5p�^�VEV��8s�: ��0��*	���ƈ�t�����e/��}�ĎOfDn�]P�D�����$T�S}��ܑ~��%�q��L~df+�o�7/'*Խ�֖Y�g�G�u���n`XP/��N��b)Sn1��,����ܝYTN%�.�刾2Kg+ٖm�l�f�PGg�MW�ġca9H��d>����2��l�#%Q%���!�\�$u���c�J0i�-*�b�
\�ڔ��0��Z!]�!O��x�0�����y�� w ��C�ቢϺ����3ԟ���+o��柧 �2�Eem"Ѐ<��gKĽ0!$=� ����?��B�7_����C�C�� Z�C���k�fȳ�d
��Ha �ku}Xkw�leq\�6�eO�Mx_%5%2���&�B�m]��\�*Eܾd��ͽ�
&��6?�N�6��xwZG[�^��!lU�����̣��cb��m�>iA��M����(��ӧj3�0j`�����!`�-=�s�����<��̊�\�K�8��%�.?m[Xf���'2�7��eR~A=F�bD���Td�w+��3�����-�+�
q ����x~ e�F/��,�V� SS�K"
�W�(k*��
��_�Ěl���,I�$�S'���Ѹ�Gހ��i}����E����$C����Y��\����K����0�|�r�Y^�{�����YW�R2D밈Ucy�A���!���/�GhS�ҽьPHQI�TF�le8��_zs�]e��H!����{�c8B`²��U<�<ÖWY&�FF�!D񎿋�I�= �����[Kuz��7a�!^8��]�%ш�}�"(A�d"%A��"�Y�`bߎ����� ��pQ�r��2z���iF��&H�^$wȚQ��d���K����Q�:� Bd��'�za�0@���L3������>��:��
!ɋP��`���!��,��zF��pG�¸���f�bp��H�g�_r�\���j�\�}��v�\lKOSIxWqsn� &�P|O��d�]�M��@�Ȋ���"j_e�g�1�:�"�O�W��
�&O\$�����Ν���W�u���&�!�z�͙��r�E���:8�RQ��d^�>T��5���Y��v�R�,Dr�'��5Ed|�O^�Xbh��m�H���~�5�^�8eS�I_�>�i�D�Cz"����_�%�%<-I�5�*R m����ai>�oy���W J���O�iޝx8g��={8��8	0�*8�/�
�>�Q�w�l?� !�;�l5W��D��pW3C�4lͩ��$ ��'�"7%����˵��Ԓ#��]Z����!��cUF �@�,�d�����8�,�s�_���V�Jף")���Ô��-h#]�v��rx6��>0$	�cQP ��9������'���[f.�đ�?����j"���<]�lcϢ���at���n5djI��s�py,�B�_&�vh�����m�/�X.��Ư٣f���X���m`wLp��ڂ_S(``�SUw �5;'r����7���G� R�X�6�|fN$4�-B�5�A"��M��Q����cFK�5�F�?��v)���u����
_���?p��7<h�O����f��f�Lػ<|1���	�� �W����c�h '��,5�c�'��c�Ø���,���>�*e���G��;��{�w �4�f�Q
Խ���L�3��,�w{a�b}ܭmξ����ֻ�`A����+��[�e=�Z���?�iqbO�ڣUy��t��X���e���71�*�WQ*��KR����\�ž%��eݖ������H
�:)0�7Uke�L�u�Kۂ����K��qӱKlj�n�j�8�'��5�7��G��'� t���
�i��sy5�)!�#^����s8W����������N���&^!>���v���=���N��	��l��P��Uz&�v�U�[���+�!������w�N�b[t�߮�JKe��ty���kVe���5.�+�փ�6ޣX�y���&j��L尽��&���Y&{��p�3�i���f��M�_�T�X^�a1�/_L	e�@���<��tTB�G�=��U[,q��I#�E7(�����H�L��5������k`��`a��mK/�K��$��;�S+F�{B$LC�5��J�"����sG�8�x�|t.����ܿ�DS��)d����϶y��!z���x8yN�g���USe���@y�3Q��| ]��>�|�� ���씑'ÿ��d��|'e�Is=�ލp	��H��Nw�����yd�}m��nZM��x
���aı��'�k8�惙/^1a!,8%�n��Rr���&׮g�Qv��	oБF��D����-��\�P\��J��P*�FC���,��L�2�J�<�A��>�\rxɘ"]�y��D?.h�T�e��ncO+;2G\�YpM�J��f�����~���n� 5~��5
��ś�t���>��S�s��i�QA5ժ� >[V1�
��t�_W�e�7�0�`�ń�n�U��3����">��q#,o]#�
��T������|�	������#J޹�!	xyv��4-]�(;/74���0�b�^o`I�{=U��Yc�i����~�����%�x��?8|sG�t�/�� k�1�i��`�f���p`"+!-�eX;uo�ǳ��Has>*^�G���`I�]�$�[;�]�Z������5� >�ޭ u�/ħDG^�Zl/�Y��;��ʻC�o�s]|/�@��)l� �ݾ�2D(%��m�_�;�wizۖ�mcsR�'T� �MrR�)?�b��@����B�'��$��:�Vݜ�J%���"��_�p�#Ȁ�O�k�����ut��,�z^�P�o���)H�}��������gV����j�
��uųq�̽ Rΰ�CD�¨��b�WH�j�)�Ob"C�RJ���a��A�1��d7��-��g+7-a�ȃ�V�"�5���7� lE�$T��><��1�-�j�����\�b��(�]����*aQ�mC������o)�GrL�?�7��P����0�CI�����(O���� �@	>x�,ts��:M�� 9�-�٦�
+8"K}�z^�K|q6L��+8���N8e)ɖ�~mU�m��74�N�* ;E���{�1e���YP� �����Y�>P��ZC&>�m3��B�����k=�t#���V���Uc@%�A΃�	���Lzp�]�kNj��>=:	q���<��9��F�ݪ�\�Hc�]?ʦ�/��wq�݄�f��0�M(��T�j6v�I�j<��,�WtO�S�������l�=� ����)E�%Z�%���b@�a2�K�ǣXs�����k��j��v��_m��n3��X�Pn��%\fR�f���FzO،!%]�������	>z�\G��<`��T��&�$@U����ͩ�Z�&%z��1dx�7jd�g�\%�S�E�#�t+��wU1R���=��Q%v�+��"�H"M�k���}�a���@1��x��
�X���B����0nY�%�3v��
v���V��_sӝ�f������U�{�?@|^��`��G,*
(�p���f�<��JW[����~:V���Jzi߸��f��O���;kT�/�ʺ�T_}z�N�#�F�Eڋ�B�_���e�������5Ҕ��Dï�*	��%��Q�Q�f��&jW��N��|O�&d2�G?a��v7̢LJ����[��d��Bl.o�ߝ�}���i��\���|֭w���Pc;��y`�C�_E'��n�2w	k)b��+c�x�L\D~q��I����Q�T��(�ҁ�OT�N�p-T"Y�^i��7
���ƥ[��3�$�Mc*�/. :U�W���A�y7]�O�3�|f�d���)>�z<V��B"��������Wm�
;L��S���y��췠��U��tQ��{e��?���/P�|��R*�E�.'gs���bb�3	!�h[��W�}�^�m2&�?���4�mu����fK@��_JU�Ժ,V��2 Ko���^-law*E��`H2,�ȝ�=)=_�\�'X����+*ķ�ϋq��&���C�A�O�
�[��O��SoĬ�I �#'�C�K?�����RvK�ƨDp��6�*(���)��K�Eb~�'LY�+>�\ ���X�Aa�x喙]�|�w�9`�9y�K�9��n�-x�,qZ}-	o�	��^)ꍧ�S�S)�L�t@��AGd�`f(K�s�b^�/7��C�g�HcH(�-�*K�잒����6�
xP��4&wmB�3���U�yc�#�&V.(�,�,1w6��Q��'�!
0S��/7fsϷ�i9��x����m.�D-Ar�#G~yؑ�pA\���Yi�@i_dw2�&H��Z|���MV���jٙ�w�r�����67�/� �R�br���� 0��RKe�r�f,}�����9��VZ��W�A����?MKQ�T�Ə'{�(��2����	�)�حF_�#�@�����r�T�G~�v�I�t��z�|^l�����r1�s���m�i� _���R�!4�I�XZc���3���Q�nJD9�E�����G4�u�m
#o۸�^,g4���<�A�ma5���Я���y�6�:���ɟ��9tV`��v){آ[7�˽$lZG�����{��:0Mp����A��g�'��^b�L�����B�X������Ui���C�WY�y���	����E-��/�/��G,^����9�|F���Db��T��u���7���Q��!?H^�%����:9H�q�n)q��.��X�j�@2M8dn�G�9����������;��Itb|c.�[���T[~��`�A�d[^�+�Y�b��J�Tʐ�Ǽ�U�pˌ�zZ�����pZ�A�����qө�n�P��Pcu=�2�
�!�P}����0[��[x��� �|@��ϓe��gHQ������?p}5Ro�d ��<<�+���S�#�ws�p�b��~(��i+߃�GE�H�0�!g��瞗�;<Ҡ!V[E';� ����^A�S��R_ׯ��Ol���)�j�����A���ߎB�>�T��r%'�ʢ	{����ڧY����ߡ��>{�B�F�����-l�<���W����冻�h��&������9N�]�8�|��J�^������=��
��%�`m����&�ww7:�9�=�����ʠ��cbp0&�#��A?e=�:4�tችB�u\����ޚ@��vkd�bd��%��d������.J�1F	�b\M�>�����rn:����d"����s�`o@���2�ɸ��e���$̓�u��.P����B'����%X��L!KJ�!Y���	6RǕ�O��m�>�R�o9q��^J#��y�q[c���+y$or<>mQ��(�8n�$����b��j[u�rm<���[���Xj�F.�����I�S]�JT�F��taJ�,-���'��N�R����t9�MΉ�y���PYaq%�7m�b����=1�N{ʍ��@�������[��񱼯�ف�s��M�{rE�@V]��*G�ۺ�{�W��:���a*l��P��E>_�!Z�{���\[�NC�Y��&�����U���Qx�-<�����7���҄~n{�m��!���߇5$�����c �^-�Sj���@�Ft���њ=!~�f�S�6��,h3��De	aa��eV�sO��b2�^�E�ց� x!ie#�m�p6~/3�0~�mO[mCNS�_:��}I��"��\o�B1��õ��?��Ls��M?l;'�d�Ǟ���q�d���oBL�O��6H�=5v�b��`����f+m,��	l�37�u
9d�`�6z �
�����r����j�9�3�	������9��Jo$�����JWN�ȅ(3��}��:c�mtY7�G�������1�Ri���7�~`P����֐�-�9%�L�g��I5,�&�}�u>�酏�ʳ#4���OJ?jJ&��7��������6��2�+����O��Y���}iW�,��H+��6����<��v�P�� U2ǫal�u��R�-�e�ӮE�e{�U�D�|,�b�.���WO?ֶ����4�)]��_�Ʋ�Y	Bh�D�"����]:�#�����E��߄�ؼٰcpg`w��3#�ѭ�,�X�6�#L�O�
d�"[I�yY�A����^2��!= 됺�������j�Ul�]�q"��Y���I�����$B�*o9��y�
+(gЦ�2d+�.Ҫ2�[Z��%E�l[��ŬP:��X��n�-��O��S��L ��W��l�&qgRY�s��0���.�f�.&�mI8��ܼjچn��)�;py3�W�n#Lロ4�ߢ��M�oh��$�C��88a�U� S�+�������E�R�����T�G�pC��4��+R!Weu.�cCɈY;����Z�4?7��ŝi0R_��ubU7	N��Y��iS�(2�`��O���E��Յ��P����:���+š���VP 5-hǳiO�)�x�0d�3'tRՊi�o"9g�����1ɞ�k��4\V�k�W=kuȭ�8X�;��4f���{��Ն�C��S��P�I:Bl�����a'�z$b\��貉[�E���I裐�ei��	3��G�A]&("��
��|U�G �+�w {�(\|#)�x��>����K���ٟ�����]#(0'��Փ;��+�G[B9�����n�z�nQX� ��F��H�^�w�m���4A��.�,�Ge��^�,>�>J�)!ns�z6���՘,��U�inl
z�my6v��K��|���?v����t#	ͶY$������P�'��}��;������c��Z���LB���ؗ��w�����{�G���%�r�����
�5W��E�(�ӽ��A��L��R
�k*4عBP�RZ�'o �����R6�o	��P���E6"##��;���M����&)5�>�,@�.fE�x�ܳY�2����}��x|6�*���i?B��"2�f�km���؃[{�,�J55�3�s��\���'ux_�'��8V�U#S�;��2?�3}i�lP̯����O�����d8��D>��!({��f�߄O<�3vPck*t_!9F�J�b����B0��q2�A�H<�&G��H� �?j�_���?jӂfG��{�>~�<�VJ?dt��x!_�*���X;������@p���%�)Vx�_n��/FB$���%�/5Xw��K'b�+o�0�=t�H�dk�y���,n��Gx;�g7���^t�%���7����eb�06t��c���P��&��|"^9ԁ�xU�O��u�k��@n�NE��*�-Dc'����<�4Q}�P���ũ�RW��/�(�Z�o7�L���o[�V����R���?w�9��C?���U�q\��;��Df��Q����;�+�2v\}ڗ��ԡv�Y��B���uQ�q�R��W\
�Mcho!�;��~W�5���ܫJ�P��y�̯/�^>�V��gmxN�t�V���PO>*!��,�d8�q��R[��ɬ+!K��)DS�w�t�WW��Kz]U�[#c����B  �