��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P�[�?.��.��l�I�2��œ��=��!?�H�xU����n�C5��ͦM�!�u1`�z
���ق7�ђ�v2A2I�~_����>U�8��sy\b%��N�i{�����9��,�َ�Q�n�mcޝeKЙ��kF���aOu�1��)�4�vV�8V'�e~�m�=&%)��}4.2�j����x�\�c+�(-P��,�"?
���fѢ<�I����}�6k��g�?��e��t;���N��PgA���V�(z�c����MUܜ꩞�~��,@81�}D "�fL�3,�b�>
ti��c����y�{�-^�ox��=K|R�cIn8$N3����9?z�.X�{�)���y���+h�%�(y�W��Dy�9��\�\E����bG,�.9�rrp#zb_���D$��y�<�T۝��ӿ�1|(��(O8�A�����u�k�u��b��K&�˿k|�,����?K�{�N�� ��[�x�#�v�|�Yp4�{��X�6.�%̒���/1{M}�q��d�o��Mܻ�w�,�������
��Y�zP�b%��cy���x73���L��J�|^�]�.0���CX��'�D[�^��8u��\(��&h�˳�̥:�U��9i��M�9����u��di��?��~\g�x�Pb����6�B�6]`�pUZ��(���p������L�%�_�ȥ��KW_���<��t�zq�ڟMi�d���0S,FNzĈ��
�T�i����2����rF���%�NL:e+C�j�2�8C+�>��SQ
�s�"f��~��lj^�?�n��<�t�`%�����{��V�n��a[�VӚ�9L/�$�08O�z�����z{�%�����A�#�i�%�0	�U���b,�D#�����(�z���F�epnv�U�� �?���a��>ŷ��)01= ���-�"9%o*8c���և^���i�~��l��>��އN�mi�oJ��K�G�3K۩D��WJ�3H������(k����/�	��2bnB< �d@�[u��47�1���Cզ���X�hi���������u)ób��k@��I�/�r"��?uyuC��J��ڊ'��:�dz��������cpY�4&~�����w��_L̃��B�`��J��&L�l���h_%s�ħU6w��xP~(���C�������׽I �:mA��u��v��v�����c����x����"H_��Jxs�G�<��e\$e���õ(ׄ���?³� ��A�]{E��<����WR���֗d&��6;d�)��p�:�g)p����#Y�����{��ڟH�ʮ%�&��.�$�͖ ����ð���JzѩD#�1�kւW��=>�m4�Q
�yAЍ�E��3�g�^F�Ztg�<�=�G���t��שP㽝�%��9.#�[�K����ݸr��7�ɻڞ�����U����Y+L�O �(��<m���)��k*��N�)����xn{��2�]�p/�+A:�ء/�E�o췟�%��l+j���cOT��j=��+�3�۫��ӮA�~3"p�))�e�)L(MdM�\)��4�)��P���	�3QN*M>P�t�����C�VI�[�I�6���"E���P��Rlqچ�x�.7Ϣ�4�Z�{�+�m+��{�;>�
��!��h�6����H���-H��rTa%��;���ͮ$"��Z-���κ"����D�s9R���f_��*a3�.}���H���:&��' �a"ׄ<ӼN�T��h�9�{(d��x����r?��y�!_�ݹ:����.ý�&f���3�Ք���ܝL(�-�h�0�0�A�k�e�OA�S�e���PPNt��v9}�>�_��~����2M�t(bmSvK轪�m�,�Y�]/.J���`zc�HNTMr��6���^���x�Z�f�`�3�x.�*ƶC�g�Kɵyȡ�*�ϓ��HI#�F��g��W�P�1�\��d�۠��%�J�ߨ�+��EM ����eQ1HS�ɰ��(ٵ��ڐ���h?�
k� ���֕{Ȱc|X�q�nI7��\����UV�	�%��!�3�	��i x�&�ߙ�a}bf�?uuV�o\q)�O �H��5C�|3[�u8]�#$�B������p�P-o�ml�1���Ab���H�{�(���i�C�	Q��V'�A��@�"E��A��V>`���o���������-�O$�$�������R㓴jbA�׸`���s�l��B�h��(��\�5������Q�����@h�WGTg#a�\ݯ�0-�P}��]��Q�X�.�xħk�Q#�C��^��x0�Usi7)��w��^�rJ�qU�ن�\~rg¿a/Uo�-���h�k'��8��_9���}�ņ�Nm��:�օ�厎�ɞ-�$	��߆B��DUJ{bsc�餮�J=���Ue�y��n}_hw /�*�<c�Ж�8p�pY=�IҚ*��z�ţ�e����"ˌG��^�F�\��lS2	��]ȧ"�J-e�����������>�αCy��T�(�I�x}���S( X���s��6V�����Q����ADu�iBj�(#�UE�������B%�RD;�*!ܣ��*gm�B+.#.�l)f��s�e��QfA�o_�lL��%�m+��W�:�����@��ꈶMo����Rl(����Z�eM����{�]���#_�i��sg��VzN�k���Y_K4�؉��-H8Z�a�Ş���X�a��RNJ��+�c��ɥ�R�qY1ɏ���E�M��2�א>AdVp����=�Ze�(�v>���=������oOӵ7�4�Ͻ���q�[�7,5��fp4(ڰ��Zo�󥂋����!��9�g|C(�xc��M�b�����6�M���,c����1V�Q԰��#w�DΞ��h'�	0���t��ΐ}��. ���3:�:I�H���現n��9q�cM�Q�ڜ�_��y��j,�O��p���f��;.�[�5"P���v0&�E">D��ߐ�F���8�h����=��,g<s��O&���s���3w䅋 �I���is��e|)�_��n^���w�i,���C�:8[`���6=����$rƷ#G"8
�{OQz�Q4
�L���Q�;
��}
y������}��L7�@$�ܿ`����p�
D|%��CŸ��ޡ�2��B`�ƭ��ֹeq	*NEf��I�Ϸ�Q1������_�ZV�x�q����Ÿ+��3��N���.Wl��N���
!��tīx�={jMt�g{����W�"��a���uk��`�q�U�: �����l�&4uE��j&�y���21�'����
����8L'o���1x����͘�̛/m�K���h��8���J2�i�.�t�u3�v*�!$p�I`���qV�d�F���̌��
��[��ܶu��V>�gHWio��]����C
q��7�/n�^g�ɚ�^ӧ��z̡��Aͮ��'��JX<���wtL�'=h����#2:i'P��T4�q2sW���xN�E��I_��[�����ڱ�?����*��"�Z�}W��#*1. �A�I�HIK1��Zc":	���͞VY�c.���*|����<=Dw8�m��,za�<����e7��:w�*��B��@�xgf�*ſ��!y3 ���%dq.�g6�xDw����0���Q��o�L����t;�ˇҭ����ڌ�������	��$Q��O�;Q��mZn؄�Pv�L�\��3�X<��H	A;�Z�^�{R�r��vq�It�/� ��_-���w�ӭ�����vo荬[�x����;�32$�A�S�GUk���ڮz��\łˉl�!uS��n�
�3��q�dٖ됋��8�{��6�D���|��ޛ�N\�
5\q��:-M)(2��+E��j-��X'K�m�惩�Ҕf�#�}��ږ:]�d>�k	�'���톉G�B-))g˙[p��AB��kp1�H<-�FɗO��*î�=}��xM̿�}��ъ�E�O���H��?!�"��2�Z�?"��ݔud��tbN�q�� a���R�\���#�	��@��S�,����wqx���(54�y�qkeė8@qk����̾��E�t�� !�o:�=����^���7�� 8�tWP�,�� �� �M��'���S�k�rG�|�����xal�i:���Z�\�����������qS��'>�N��s�
����&�o%����a�Eg������_�#�7�W�c��>U��V���A�Q\ïA>���D��Rr����?��E{NEQ�nԮ<5��l��[RJ�]���|��e�a(����J$���U�6���a�P�`;�>T@��3�Nv̑�_��w�̹k�����bXң#rc^K�"S��.B���R��k4�ƀ*D:@Tηh1��F���}�� ��A'L^��3Y��.��	�8�u���.��g����'Q�k�ٖ÷+Ƥ*�)�7�WC*�q�s<�n{3�V�\fݒ��n�ʽ�	�ۋ_i�k�WBҟ���=Ǒ#[lI�;�$��Ꜿ/�����m���s����Tr�
i��W���$<Ѣ�_��k��2���.���P=k/3���}!��6��=�\��xD�ww@�21�,��d�G���h���n����Uiˍe��c�E\j�W��Pz�K���Iʁd�)jޒp �M�� �(	�y�P�T��	�[v��ď�`���2KՁ�����`DC<*���|o��?Q�/\Osn�P�M'2��v �+�(x��0N���
{�E�pM7�W��R
nP�ַ~�\���,,�F�B���5�qNl����G|P�|w�{�1ǩ4w��,%�l�q��-�}˄X{z���U��=�*y�43�g������J���Q��)�	/�)vp�5"�V"�!���0��䐥x'r�7���N��5���m���O{�(����<��.����n�V���ĮY)'�cF���C�Vzw�m~nC���"ߵ���P"U0b��O���Z�Z<���}���q��XJӗ��5��Tf�����@LGRi4�#�}I�8���:���u!�`�4��2�T�.���N\��3~�)d������K�j��-?�������(&W�;��ۻцB�L3�ji�)ʥ�����G2)P�}�4`�g�vߚ9:,wR�e.
�&��䥉P�$���r�\�棇�g�u3�Z7Os~�O,Jă��5��6���6qt��)��Yh|"q-�s4�D�>�F�æ�MA��4\h�<�X'����y|5<�M�1-�+n$����=�9�}����}B*�Ip�	�~���b���8+��M�L�4=����Ei^)���{���Ϗh^nf���a��:=�����q�27��ji.E�~I��Z�v�?,鴁{��Q��SD)kəCBPm����WB���N�M�Z&	+��e���j���3ވ0�EW��s*�>�	7_�CX�)�	˭gp�a�M���?Y�e���f�֪�QB��&�UYQ3$U�������V��J��BwdF'�֢8ш��6�`p�lE�+X3���<#2o��:����H1��q
Wq��y�F<�H��L�fB���v���g��6N@���G�*{���uOȮ�v|��&&�F����a�����~����w�6���� �}0�*g�� W|iߑA)��������r�w ވ�׆��'Z����U��"�t��N������0���.�� Y�M�Yi�bӓ��,I��l8hj����+u9s׆�QCm��)r�e���q�v�	~F�W ."0��5_;�N8��8FLJ�ģ�<�{�]�aZ���.��G���u�u�Y�A����w��()��ˆ@p�78{b���!j��"U��U����e�`0��X�ۯͯ�lrU�I!������*��BqfLHQ�Ww0a��:�.J�A�6�d���N�촪�=>�M�>�.v�2�s2�j�dח��~f����'�4'@���9��SMt���c!����g���G�y��'(�j��ا6AZh_w�nVF4�-�hNE���M�$�Ɖ����}���@�7Uwl�RIN� �.�$zXB�\>b���d*&� J�zǱ��؁z�櫖eI���z5��*ؽ�i:�J	"�2���ѵ�xES� �Hb������3��_e����DϽ�23/сc�7!})C/L۽�g��-J5��aE�ԄvG��m��T�\��<�������`\J��#�U����޾نv��W"�V���:����":Fk���b�f�DeWVxӋ� �)Y�8%#�Xꬤ�%�]�^��;��jl��FMo|)"yY��6�}T{��*�9�,A�Vs��K��J_��$	�Oب��-Ӌ�Y7�Q�)�\�梡�L]mP��9<�˒:��;�k!7*�y�x�v/�(I o�J?�]Z{��M�C�u�"n$��<f�/�K.��]�
�~���I'6o		M��:99?���2~� ��J%P�Pq�5l��N���mz8$�H�@\��Y������χ[0���H�W�-�jqwG��0-&+Bɇ }�l�1�`t	Y<��*�'�����ӗOeV9SJ���x���H���gn�r ��Ң��D5��
�b3���^�8�� �Yh�*�͠�����7��3��k髁t����.w&�]@�Is�I���Ɲex>"��X�ʐP�5#�%�������`���2^�-�L�!�5^����h��=��?�y�&Fx�R��e����W&�W�RC$s�)��xY��S�S��/v|��
�r�-t=�5v�1P5J��|�'��h������ͬ��R���x�e%�+2_6$J����pl��@0�A�G�"�[��Հ�����/����ȳ���%��i��{$`��p�?5�#5f~�-��_4�]\��*��^�v�G�����v+�~�����{���6�ƅ��:��ȁ=���@�Wۗ$$-uƻ�+�h����J�%������a�����R(Gp����j
Ѣ8h��Xо��HfA����V�g�M�G2

�D(�|E��o@N��rg�釽�^H�<#�"-�O�e�V�?d-�9����V�b����+i$��vJ�5Yc�o�Z=i�sr��[W��B	SS9�����F�x��%r_[�����	�Q{�Z ��(����K+���L�t�i)��9_O��B�jgc�
��܄�=����R�P��1�4�A� 0����VV�� �&���T��۰�N)���ؗ�gw�X�|�u��8B�6�B!t뤧*K�R�|1M�1���4�iXR��]���(
"k��L�1\����8�g؊�f�_��w)�\�ٓg�hZ0y�*� �fjJ��cNB6���)΋m�@T��B������t������2(�����7?�[l�Y�-�D7�Vm8ڃ���������m�$,�9ҷ@D~UＥ�=�;�iXE֤晧�TC�4��P��D���)EgNL?�<���c���B4а�`��E�iw�ҡd�J߄�q01���-��$IG�,����&t  E��ώ���!����y�۬�t+jc�E�'0����26��PP痀�;O�T+��1{�˸�2�� j^1��]�pK�_<���`�=��4�W�O �8�N���I�������U�,Pa�j
j!Kfvre��!�x��s��A� ��*�����֠�3 �Ju�\PZ��reM�D��K�i��ƥ�<�z͘�L������t�B���qH"�Y�C^�s��t�4X��v<1p�Vj�r���b�kU1�WL��dyo��� ���У1��[�4j4L:z̴��L�\�	�$
����j�憔����e<�?��p�X}�H���,xV$��z"�8��)�}�[�C�����D`�ɋ+Vedӎ��/cO��
;A>�. ��U�.�0Q� ���H�TՀ������L�w��i��s�3�͊�D3=��E
���!�1O�Z�R;��ll���V��Fx-�����ѯ���x�w�Y�{F^2�
��P��WH*-y=w���yɍyE�7��B�"����8
��|s-^�<�Ό7ꇈ�IS���������nZ5�e�>b�'��az\7G"��3]>�$}��|�����?���D(�ZОRز�Js~1�v�`S�,��5KK��B��`�m4�<ւ�N"XB	���x����J.f7����X�{ ��K�\�	��o�.�S*Kђ1��͹Fx���p{�Y/ݥ:Zj%7t���V���G�������<����Y���R	�����/PG��>��a��E�m��C��/���g��|�^B8��d�(�0�1��L�'d0�G:��!I� jmI�7�JQ�CCVOm*	)�E
�y�qz��7��LBP�H�뱰M����	BCꔐ��4���}!��/���d�y.�W��;�����tez���@�9�ҍȀ;fg8�Q=D;A���O����&F�b�L6�����B�<��H�J���B��Z�!S��A8Q���ɴ�S��f����HR9 f��=[,#�#za����_I�՜���v�X0|��>����s=J�:�x0��&�� k ��2�iU-�o":n��}:�k�8���[,��U)T�C���q�v�-;�o=*��s�3��{O��MB���%U6�ح�\ȏO~����������#%O5��FR��K�e$���hm<�ûB j-�WG�,��)h>��6v%��ʧ�}�6Oz��!�>�g��0���8Ļr6Vk��
��C�!�GaB��֞����^�쀫����4o�hE%�N��U��
�5��~����ᖧ�s��3{�Ⲅ�� ��l�Ü)я�;_�:���:������0h!2s)M@�BִuH���!~V�&����c� !�댠���ڄ��H"��A�	R���bA��#u�����k���gL�;cg��q wk��N���5_�����=�	�U_��2�T�PA�4�z��2s�v������	A�~��l;r�L�k~4j�T�L>o"J�����mm�ג�/8��6a��HR*'@�tA�]r��r?i��-"���*��q��-!`vd�]PC]v D7Z:���;���$�{��J:?��G��HE�8Ԟ�}+���O�S��'�$������W�@��q=;��������﷫�9�z����CSb��H�ԥ�*SZ���p[���N�0��!�7�93��?:PwG���\f�mM<"���K���-���<�V��MJ�$�>hO��ݙ{`=�|$6rw�����`��ơ���� �.<��8V]}i9�6{�Yr�.���+1�����<�����	���a�s%�"CY��}�(�l����F�;픥��"<��k�ԝI���.z1d�"h��1�W�d?1��� Y��wRZC��U5�G�è' �%l�:����7�iʑ��6g�gƈ�Q]�_�g�`w�t�.+����N@�/4��g�].��2�A�vrz��L��"��J2.��Sj9�켿��2�
��
�0�ɟ[.���	�y����{��1l�og=7�|����CM�q�Hh�9�h<+��Q�����ƻ?�O)��V�~.aQqRv�V Z���·]�o#$?�C��X��f�-P�Dy�p��b5ލ�O����z�{�nyD� ��q�cJ��8\�j��W��jY��u�o�~Ƙ�N[Ƒ�������p��l���(��
t[�_vkͮk�I)k壘P����{�n*�h�6��)i�r����Z��g��@���z|ad��Gȱ@����~����4�H��_q/�'ck�@/�;?!��zB�z'��o)��p�Пj�pLN�``#������"�v�Mcp��p�Óf8��+���B�(��2��oH�%�̜����%���4 ��.��q.�ʖw�l�H�Z,�ͥ��}����;�F���~�P+�͔;ĭl�R���W_�m*�AI����$����؅-��M>�XB�N�c�Ć��W�u���#�2�$k����i�7�6�'L�ll�@A�ͣZ��(
^�~^�����"�e �
u�̤J�)M,�pԡi!qc邾+�ti�ԟ-f.��t�J]�5���(��(��{z��[s���s��*R1����ފ���	[�o�d��ҴJ�Y���w�?�j^&4%�x�'����Hd� "W��;�֫����:5y��Q>��n��{KY<������PΨ.�g�����z�Y�۱J����ԣF��K#�+X�0NTa��6�����X~fO��[Z�M�h6"Fwj���WHo��H�9����o++>㟔	�g4���#����}jI�M]d�)��c@�|�	G�%�r�i���;�ڱ���B|��8��[��E2�(_!�!���.Q��<3�g�	��Y�.�.�o7�ρ!?l�,�S�P��ݏW�4A���M��Z�>���f�9_��)H�@������ �#����eI�~g�"Zc/��Wʬ�ޅ�4h�?p{K)v2�mv���
2)Uev��Y���ח��������`"D���}��[���H¡T���8��A��2`g�k�aIl6��N=������!{�Э\��g:�\���ݒ�Zx�mWG_�Tި*�ן_G��~��)� �����������M��*O���s��r/��A1�#_��n��\��d �6?f��>hU���[���8��P��'u�/^��d���G�,46���PǇlb���B|���f�i��k��(�1�53(�*mh5��?#J�æ6h����'�}Ű�n�`}��<=�-�"����&��߀���P�f�f>=�|n����N�s���^+s���tyZ�����"Ԛ�]ßO?,!�i���<?q=@X�gxֺG}`���I���o��ȋ��u��p Y��,_��uq��+�.�]����|��Ub�/�ܶN/4��1�l�6�)�_dM�j���y��p���x�(`ƨ�[��JV�$Y�O辪�G��~'����P���N��pgOzIv$�TgYJ�Y5�0H:N6>�O�p����Co��r"�+�m!� ��~!�>����]#7W$�z�u�R>��ȝ7y�4��>�/-�9�f��>m���#�v���*�G`	�ɧvk��+_�Է����ѿM�`_��r�xu��S�Q���2������=_M��h�U����j�ԍ���<��;2F��"�pҭsW��C�+�<z| ��8>3}���,�#
�3*��SP_1�j:B �B9�/�ri����'~��1�@ы�Gh����=�{[��0�u�`�_��@��>d���fJ��#_?�g�,m�a6H� β��|C�oy3ݷ�$F��L�Q��d�P�Z�h+� �(n��l�vYW�wz�F�4qSJ<Oãk�M�,8���Ǐ{Ck�o��Cֶ�+G�KR�`����{^��pM-������`��@Y�7w2U�SB^��G�~l��K�\�(�ɺ�p����KN�~��@����T1���=�a��ėi��V�ƑA�*6T���2>; �ÑY�Kf\�G��q��D%�Ƚ�N#��T��%F�1��Oehb$Π"B�������m���n9��A ���@ӿ���6� 8u+��Rw�v13H�@�S�	���4jwS��q��T��$r(�zN��+�G@�ԟw5��Xp#�O��8�e���GX`� � h ����^vKL�f�³5�0�4����S��IzU����˭���<��Z��<8�E���zsu����0�!��(�.��9��.~��HT��s)[-U�x��W�Ѕ}]j����/ݺ��Ǟ�E�Z]�ڠi�Zzg�o�lc���J�N�{#j��]��z�d��L�$w|P���/�����Ԩ��6֮�9�B)
FϿ���k���!K˦4�a��t�\��r2d��j��B��S�%eqL���9��s���*̏�B�X���2���:�O�&�0���n��n#
w���あ�WD- �k%��ı��~S<�������j��d0���<�kΉ�p�p++xL���Q�%+É	- �@3H;�ah3���'A��,� �02R�M!&H�H��`�������Y#���OB��,���	61-(�zz8���jD�{nPF"��[��T��.̼(w�c�$ҳ=f�ޒa)v�����xl�+5|�g�	�=�Q��UC�D�M�:�~04w�>�i�._H�8B�k4H��aVǇ�,�i%7�Bj�����Q��ȕA^.��{���*���7[����#N��IN	�R�rY�\#�5�M4�ș������E� �TL���-�n��7�g��KqT�ے�Q��8��*��u+� ��:�����w��oY&;�XzRI^e��[�����q�����m8W�cr���ֳB��B��@��c�����
^EN	&�[Uc�tF�3t%�E-rI�E�eKg0�ɖ��i�l<̒܊�,��z��L@�z�,�`���,aw��� &J܏0(�xp��O�1V��W�. n�����Y�&�*C���N��M�ς�?���?��A@?�l�!�|u[�/nč=�K�ĩ��n���h-M(t�Ե�9}���ZE%�G=����j|!2�sx�V�.V���z]�]y6X��4
q0�6�����c!�O�4aq�͐��毕��j��/��*�/�(�H$')z&q}j`rv�e�P:M�y��3{X���h� '5��[%Z���G�|7��[HgYx�gcm��&߈|`�}1��//�����:����5�q�-�c����:�sK+q��]��k$3]c��v�,�j���I;��I��ۯ�ǁ^�SVKv�O���JȀe�-S��|g��i7���3j��Ӌϴ\�Wfd}�,�C��73.��sUx�g�������կ�t,�WW*V�h��p�[���	����HOǆ��"�#(c�ȿ���;N��
E�
�WX
�Gq	 OȦH�m�@}�1 ���J�c���Y�s	�2N���F��R�lP��Z�ҋ�[��e�N�`P�R�X1c��#k���U^�#�ha�De$k�$��F��]���ճ��|/���"8�+� ��FEJj��)�d#�� �Se"�k%��ⲽ�o2	�C��tHu]�2�\�$ă/��]S��1""	�BāF~�=/�$�� 1k,�c����Vf�>q0
�&o���c&�LK}����n��FZ�?����lFT������c�)�hUgOگ���^��wz�u��}7��W������e�D*���q^����J�IK�m�&�
;��;�7�_�
	=�?��[��(��yܠ�O���+)UZ�C��E�]X����oaZ'�zmA� xˏ�R�=��{;`v���&�a�� �A����DOpB�����X�t!�zPKtTG�߇�0�X��b�{�f���AQi�H�jIp��p�g��"�s�F��>�l���4�S|������O��ϳ��"�cF�6���M~�=JՒi[X�����L�� � �n��DQLv���d��uG�W�@m������"�E��69�e�h6	�FU1[�ڎ_��0=E$�,uDc>,W��c^ +��J�њ^c�I��dH�u�yf&�LG�K��d�ݨnq�t'V�r���V�a��r_-@H�ҊQ1��LukB�ʴ�0��]]���)�^{�f7|�ts���^_t9O$"=�¬��v��uX3h�t2�3O~>�T��뒝]8M�DE>������i5;�٭b����u��
[��h� �^@�Ь�l2�����adKڼ#`�>�2�"6��>�u� 0'g��S<�N�<f�6�*tjk�M�2�'oV����6�Jr)��8���8]8�ݻҽ��[�M��O�4.��4@Y���c($�]+ѝn��CZ*�A�"1.C���c�dn+8�.�4��ϸ���6����ٽ:��>���5Z#:���Vx�dj�n��q\qdF�Ƅ5�Et�@Fq��)�)��-~w\��B�%�'�QK�����c��,���f+U����g��ܩ�	���ʴPE�Q���p)�gkb�kKQ���f\��"��U��Ra����s��`����:?{���PT��mh�#8n����O�J���D���񗮀S�C
�\-%��H6y���L�#	�Gёt�<���������X�9e1r�&�@X����nk�Ȧ#����hu _��.��._Q���	ǹ򷴇�Ӊp�9N;�؏&ܛ���C�~�	AڌMf��85�<@�=ZR�X��QȽ��a�
��0�b񝨔��V��;1PQ��8aNc�F�6ѝl��íz�OL����$NAF{�"�6���UJ0q��!�p��"��R�p��B�v���P���J�P(�9É%%Q�ګI�Sx�De�QH�Q��_�O�ƽ�k$�7h��8�G�}�E���O���I>x��pݔ�t��%�R9��+��~�d���;�$�(�vͶ[�G-�������ɿ�R�?�ɡ��Hm|���au�s8�
�?�{�dβ���T@-#A�^��(?[� ?(�8���(#��z�@�x�wP���{�L��h.b��R�?��ty\�D�:/�(S^�4���3�i�ꔅ������#.G������#�N�$R:��ͫ�p���VRj�ϝ�=���WMH�7�zW�iW�D>�/<ā�A�PT�B{��&.%�=��FΆ"�T �t�,?G���GT���v>`�jQ�A:	�NPY(���}�>�H+�Ț��H���������\R�{q��nl �V�/x���~[u�Y�z�\3�B�J\=�Ҫ�O]Q�{?@ӤK�K�����fA}*c�|b'"�a���mL�7s�"���__*i�ŧr&(,��e��=�k�YZc`j�V�j⹽�ݱ����� A�V�{�̠I���&C�}�S;�V�[i�+(]�A:{ѐ����M������e:�	F7��q��T�F�o�6��P��5����n|�˃:C^�7ߜ`�N��A��ǲ��ױN7{�8F�}��:�P��k�c���goHS��i6v�g%c����&x�BxڪqW��u�yA}� s�R��������+~�`,�m&���!�� -�"�l���r=(ϔ�����^�̠&=���L�)��<z�M�L���̊��cy�,���ۋ8����	Ů�!#�V���X��9K,,��8nu�Z/�4�nB�)�4ht�YY�:�	[���A�uoAd�^��K�J�TUȼV��5c)��2ao���Y�j���Ygon����������s���(�`��������X�vg�u��P��w�%��`���F	�i��G�q��լݍ�/��{ge���a��&�d���=i¤A�<*%�?F?�V?���7��U���Nk�U0I�cmE#�v{	�&����t4�LF7���"W1��q�(��f՗������ ��Fh�����\���Pk�r����ܲld:�g��F���(;-�=�]l3<���Jǭz�<&�ʐY,*��Ät�Z"�Q�-c�=(%�#��\�����9Va�ԍ`F&i�m�膎G(\-P�^DsV�6�Ɨ����!��O����гL΢�����Ő ��J�@�a+`�R���
����Pp9�ba?N���c�0<)�*p�GmԞh�tW�<�6��Lq3���ۛͧ��B5(LG��a���̴�j�2h9�y9�� �w���N!�y���#�j��(�
�\7��덑�g�K����eS��_�	R!����;�t1	�=��B�ـ�I��G.8t��*h߹��^u����Egc8��799�(E���[��>�ϵaGte�Ο^u��V�@h�Bj=o�[c�#ň�t�W����¦�-f�;;��n	��2$���	#x6�\i:��w� ����B'Պ�d�$K�h\��%�u�Z��l�;EϨ�)e���ى��")\���n$��+%YT��iM�9o9��J�O���qu�+���U�K�%�	E���W�D7�	֊_�|{��y|1�$Qd��,0��4�P��v��5�CBէ�*�Gu긮l��v����ǒ�mS�m�ad1ѭo���(��K�����o��R�b�s�π{�胹\(��S�F>+��{r�ץg�R|�r�hXOu�8÷y`�9�� ��L�9/�G����I\�j&���?F�xz�I*�j*nՉ�IE�!�n����I�6
����\�O ��hհu;�����d�K��iŌER��X�[�>�2���\^J�?hQ���,W���$�H)���Mס<Q^X��Q2YL*T-ө��x���=|%.�<�Y�K�&�nL��(���Q�/�(P�$&pU��Xar�M8Z�eM�Ba�Dt ƥ[¤�m0dbv��hv#rpx4���b�d<*uʋ���A�S1�g}Q$$���+1�Z��<y"���5F�â��0���խ�ff��Ұ����{ͷJ������}Þ#�'&�ޭi�&�õ!V��]_IRP2�.f��l���<�jB���;����V��W�4W�*�98�bk���7�ۢ��-��n���=@S�j��*2W��T����p��Y�Bê��0a�Ӵ�zd5bm�v�Ƒf�5���7���S�����yg��Ԏe����i(��o ��L:�J� �#q�q�c|�#f�,�.i�603��Dn5����Q/�����i���k�f��Wv3V����H�c+}Ii�g����By@p���a�}X��y��l8W�����(��JNYSKiZ�mX�I4�=*[��<�Id��vò:��v�u���$�^�:g�WO�#ꜥ]F����V۴���(�u��ߗK`�n+�� #	��8�����bW�t�:�\(�A��/[��ލ��>��|<T,����h
��d�j�92�R����@�G82}?��5��/����Te���9�J�i�Cc��XǦt��ÌK+��)�����e�U˩���_��D�%�{@��u��]9���ـ�����~�ZU�h�4,Y�B(��n����=��U�X5S75kF��:�r��7b���w��'1b�r�2!@�I�sfG@G1�]���b��D��_�ݰ�x�
��6�-E�?`;e�d�?��O�f�5P�w������;�l�/r��@J�����E��������_k0\�D�%i�>��M)Ḏ�X���$��J��&��Dw"�gj��؟�`Qs,O��$E���E{t �қ���Bcl�p�����#�j�+�s,%�N9��Wx��;N>o9Y;#�t��k"%�^kY޹f�j�����6�]�3����?���/`Bg��D�-�؈c��;�6zn���R;��Oǭ엠���� ����������O�)���*��u����*Bƽ�!Ms��΃���Ȋ�>&*��osf��ˬ���`E�_�ԁd������c��X<�j0Ty=~U/)�M*�%���u[{>(4���N}��X�G|�^&��٩��US�аb7q��־O�k�����z�'`���~=����wa٣Uzw���P�.���BJ8��߬�4~�r�7�ܔ���h�Y<L�j3���脈`�|�i�UX�_ ~xN����oz�[K�m+���܇0��sIf��I>ߩƒg�(�0��O���8݇��3M"F��іa��õߝ�^���M��!���C����E��Hóg��;�ċ_��
��m�?z0�C3�_�$&ǀS�I,U���g$Æ�Qv�Dzi�����!�}��Z�Flh���Q��=:C��e%���Qc]~�]�E��opS�X4=�uQ�x��#n����uiu�=:ȹ�+LeU�=*?D�� �D0�YT�V`���7�t��J���2D�SN��H�Ý��<������o��Q�ӯQM��7riĝѐd�N��ػ��hv"��3P%Q�7xH�eֶ�ͪ���gu-�[�u�A \ځ�ts@�M)�v�����Й+|�"f%���+�4,p�[�r�U�Xt��o��,SQ"��i��Q@=��E'!\_�0Uz� ��d�Y��A~����I�{ �@��'�ЖݓT����@�����Z�hW>�����.}��m-3
:O^fi�����G��X�p�0t��G}dV�LN���
e����^��==�,
�^�����CyB6'��B� �ǎK<q���|�t���[��Dlq�w�јYɅXBd�zެ0;Q]R8^�`�*�c���jB��%��=�62r�P΀�bRP�gzjOY �Q�� ɤPj���U:M�L��ҵ4(�[��u�p��(ԡ6+MP�r����_�8������uS�d��N�1���)~N��z�UDZ�-&�1Ax�_.�jR�RK�v�J['�=��36'ۼ�-��X)�`�q*�;��%�ʺ��w�}1�i�HQUM�qi� ��f��NH��.���U"�蛞�|��
�(�-�+���Ta�gYI�BN<N���7ֺE��&�wV]�Zj5u+�L�g�Ҳ�`�4ei������RL�������{oG��13kR<����Λ�(����p�w�ImǴ'VT�xXv~�E�:QD��� C���{"����VA:�2�G���(?^=�#L=rS�B3x�N��)��oq:9��En����a@0�B�%/�b���bg �ɬ1�eL9����,��=��";�_���=�whA��@J�s��
���I"J��o1?�'�K���Y�N���Aj�E�Ihyz��F�=�J����L���^��	ֿ󶠢�<�0���Z�ލA�؄S�����]��+��āa�ۺ�9`y{��0�&��/ʟk:���T"�R��U��_�&�\�	Qh�Q�*^x�T?ݾA6�ttMGd��v��"z���"F������7�0	#b�.riB��&c��Y?�5?�U	"��~
��1����;�]ژ�x��w�e�k���r(�i������n`8X'ߏ�hV�KL����QF�n����ti�^U+3���U�3�z��'���	}�m�@Ͷũ���# Y���W?s�$#�D}y5i��< �{�2ֆ�q�E�)b�_� uGp�����Hlh�w ���,�
��N"�\���THp�~tڟvj]�d�����5(�c��jک�D�- ��x�)蓰F�PzJ�h�(��"q��c���b�w���[_�s���?w�����'�~��Ay�oB ;�)w���6��?3���2,��Zb�����C&,��K�}EB�hT�(dғ'��Q���SN�b�ϧ��7�m)e;���aƼox	�`,��g�2������߮3�A"�XT�y%�1˓�8Q8H1%N0�L�8ŉ�F�ec;�Ieb��˜�
��Rp�@�Hm��7D���\� +�o�~S+{�* ����Y(%1g�$@��l��k(�,bilN�� |��yV��Ju+U��:׆�=$i�\�L%��V�pc�!S����h��
�b^sP�'�h�!q8q�����>&K��4�4t��#J���HO��?Vy��X�����j�B���}�Zj�Bײ�� T��R��=���"�m�	.2������#\>���_��F���s��04Y�`��n�F�
�C�����\n&��\���j;��'��G :;��V�J�qBV�[���D����S�����$P9I� �]���5�o�*^'��=���6��b��%ɡ�c�e0�&ɱF���(6	��rNf*�0��7 wܡ�V�f	q^w�C�|(�-K �Q�'X��p�c-^���"��D!Mq����O�r���~�b�fj`�z5P�b�)�����a��ov彤��5ap�;r��Y�eCf��g�[~=z��O.[�לj���z���62���4f��泳����m��B�(y��@2�i�p��hc+�?�Hq)S����:T.�*%;�-���̆s�=�;���v��i�����tLN*U�Nj�f�/{;^���9�@���FqC�2����)�j,������6��}C�uk)c��ڰGw�1M[�w:�s�׸~V-��r
ކg�u�.!�	,bR�W��M��V{P�t�7w�՜6�{�-��DK�5_S�� Z8�D����o�(��0����~�u�}�LyV����Ynؘ)(v�gHA����5ϛ"��l��q=�<bs�=w����d�;|�$����ݏU^��s��j���َ4��[���$u��Or���X`�jPi�t�Ŀ��hw�FS�����Bfݷ����Q:G�"�'H�o� ���>���2��q�^#��d#��"ivx�m5Lq��VerC�m�����p�����!D'�$���"�U�G(@�m��mL{�k�
*�ۑU��TR��HD[|�n��_�o�7HX#H�XR���$�x�ȕ�hN�A�5�߲)��"���ؒ#��䯺�e��\ͥ�.5h�e��w�+�K(nUz���t�{ujQH�U����"қ*����IC�=�*�x
U�6Sh�B��D��l4�c"ط���T�67�w��G;�N�{x�0� z�mpb��~��i�-g���!�����w�>X��ȉS9>�h)j�Ÿ���B��q1�N}\�vp���2�=\Ü��RU�?����r��W�`���� T�� � ��T�����#�	L�^Yw �L���e����K�{���<	�O�èIc����DGm��S�X{.�q�K�ƃ�;���w�9�h����L�8 �GY���0�AQ�UC�Dl\�+��l�6{�k���9���=7OɬJ�K.53���Z����ѹtL�!�{�=���%�u+[���/�t�K;�}����b=���	�ʏ�v�&c�dO@�[h�t{�������?�����`q�c��`��\5Ѓ�3�/-΍����ק$|	���K��n�?{�~�K�� ┶d�C�e����	�v�P�]+s/�i� sκ��O	\��h>��`���K�C�C�*�����h��m��7&��.�����!�O���?�;G�3{d9--e���,̴nDg���H(�e�L}3!ߜL�֜�Z���T�ھ=p�@]U(��k?�N�ZrgE��ۆ��W�
=�C��Y�*�{��<`�c����
&��T�Z�\��w�I��]0ڢSf�~0q@6��N4�q��b��6�s$�X���e�d��DW�=����^ضsvS'��"�j{F�߬��y���(���n�/|��R��G�Y@p�g�Cb������"�b�!��a[�WDh��Iz�$�]�ƀuT~�����`�B�-/`��D��+8��<y��^0&|��,�m�Qd6[8�gYzs��B�M1nP�D@���O����r��2�l"�ڋ� �O�l(�sSN�$yG��J�O�����G������Wkv����ޅ��7�/׭���.M����]���~�*��b����x�t����pD�
�V�S���.Q��O55P���<�$���Y��[��]Q�q��NS
E�y����1a.-8댛H�fa="��'V�����#�^r��gA���d�I`D�%��8���!��H��Z.| �
S�m�Q̑��k	����^K ��Ƚ���c�GIț`M}�Q��L#kJ�\ɜ�Dj�I���L;�=��� ����>|�^XT���~���
9���ቫ��B�Z���~�Um��	!�70p'�7��j{0.A/>�1g��=���J�2>�.�����#����q\P{��~���0������Q:�� �[6Ri܉ɆSZ
�t��,�����|p��1f}�u�1-q����ъU�� ���x`� n�S7���l,�p�J]g����;Wū������%�@6򔊹*���xx���qj�I@w�1{����M�w#fTk�a�������`Eާ�Z4?��E�8{kVh��:�]�i��?��A���9d��`W�Ɏ��H^{j�{l8 �L��q��&�ƃsl�Q������b���;*���Y���d��]ws�
�˿�ܢ![ݼ��.�_��ZT��n1�/�rLI}�mI iwS�g�;��x��80�>^5��<�i� N� ��yӐ�Ū�Ǎ>V�c������/]�y�K=Jf t��������ߢ�2�o8ńq�mr��Q@b�Z��{:h�i�g����S�]ͪ�0*�H��Lܓ�$��/��� 	�h���4%�K�r� snf����R��X���6Ym�>�����-:˼��2r<o@�A�q0^\r������A1�)	��z���	l�?��ç2�K�_L�w*��p�4���E���F�U�b�-#o��k�,['4�_Li�\�+�Ζ�����k��cg�h�-���
�	^�FS��E.���F�uPL�GH�����g���Ʉ_D���0�uu�ؙ�J|;N� �u��������ew��D�\3��@��T㦽���hǦi6[��
��!S5R���F����[�#��gd���æ�E��b��(
F��>Ye�O�5zȑ�C�%,C����<��l��>�P	�Ԃ�!�hݳ��u�|��xK��fQ�f��9����`ie3��U�0��{%g�,R�sHB��  U����h�$#�x�����!	d��I���|��������.q�S$��&W�I���%�C_�Ц(��f�^�(��T{Zσ��^�d<�����L�JN�X��! F"����ȼ.���i�4w��s3���ze�[-)Ŝ�~���$��O�*cC-��m�����:�֔�����ԏ"6q|�e5�t�sl�8˅Z}ȹ�����I�xM�h�����嬎�<�×_�6)؍�v��s�䇟��pGD
��Q�ݐ1mk���.��̓�rœ��N��&.�M��b�xT���b����<�P~���l�?��/:@�u|���|�%� ! �]�;�ָ��nٶ��=:le��{19V9M�t!o<��r:�S�%)��x���ʘaƮ�kU�x�	�yd^�"k�*pqَb}��RU�J
U���.�v�G�D	����)�,��1��N>�M�k�<+��>s
a��Å��� ����(kp��$�y&���ٰ�� ��RAœ`����/nSR����\�gq1-��j�����ܳ��}�9ܷb�a6]]i�á��t�#!���k�r�:�&�J�kAW����U��$�����J���:�D����{|"�3?(������}�BG���
���Hy��򪐠ty��8��uU���5z^����`���h��w�7�T㖛VN�J$�(�Y��nl��}�Y�]��b��� ,Js�Bv�������갥�wr��Q@[ ��䱎�u�"�3J2,�,$��� �­1��z�3f�E�\�F�����2��㞈Nh�2��D��7�nx�U���?A�~cr��14�aA��7W!�� f�o)n?kg7*�.	�l���O�@4��&���g�@���D_7@R
U�?�����+'�*L�,`���ؾ^�b�N
��
R�֭��s=&�94�d��_"���[w=0�pG�ku��z�6��E������6i~��y}go��w�=��	뜊�^�f֍5l���
i)x�]}^T��V�̎5Z�r�8�ˤ���`�(�������@�՚
U�r��"od7s׮�f�ބ��gw�DTA�u��YD�N��//��|l�8�@lR�]T߈%����7p����5�m/������bq�.�\��l"��K�Y�O�Hŋ�d����7�~�*<N1�x�c��ꘫI=Yl���պ���O�\2�G������\c����!���܈tD�ͼ�����P�y4sw�@k����:�r��7�8�-�,��,:��O0���mk�y��/p�9a"��h�Yօ���h1� ���Q�d%<�9p8 SP6(͂$$'m�#;��V1�pR �7�!������?�"\>���"�D���&I�͟�x슀3M0�e樚�O�i�_O
�JO杢vn�q�r�4�\È'�i��Y9���mQ����L{y<3�M�{Ww��;ԇ)G;��R���Ƽf�(pз��s+ڏi�ֽ�
�c8�_�{N���)��)��3�࢛������ٝ~9��L_�3߻qϊڼB|�C�H�G�q�QLeo�|��t�^n{�hie@���Q��<B"M�牱d�#�fi��Pn�j��^�(4�e<�P�pu眝P]x�{�^;�	ڡ$���PK��]F�g�.	�%���Qw�(��J�v�F}g��,��=tb�M������!T�\,�����a���]���:�:������8B���~썼?�y�hj4w��馬S�0�?�x!�\����󷔔_���ƫ���j 	�u��>lH[��|�* L�z��s� F�P��U�M
����제'ᑰs?����� I\V�<��%�,o��"ć���F�Kl�A����M����%=��a��H��~���@xa�hd4sɀ&�x�as!�P2�0w���|fx���-C��4o�`Բ��p5a?M<`��o���i�����[@J�-�lCac,�J�,|e��~Yxz̗���ɪ�uy�#}�,� �[Jj�L/���p��$���4��&���Y�eL"�0�$���ࡺ�'.n9�,��x�MS��]v�h"�Jl�Jv�����'R
SU84�YQ��)}�_M��gr�gC�IHs�]�>8v�y�;�q����>��	]��YK��{��BjF7s��[ơz�8�z���:��sh��}��U��4��k�^V�IYO��8���_�~��h[{�=�5�g�"x����e�粆��f}6D�J �3,r��'B�Z�?���UH��\ı�6��,�]��񦷼�V�k�󧠮��.Q�����XO��B�e�Ԕ'��;��[c�S�ͽ�zo? ���u�=�8�ȩ�3�fk�Q�1�<!��Mp!�D��(,͇�O����Ws�-�M�S�̻���44*]�/̆���|�!Z�VwE}�v���v�1�M���X���KDN��_&:dY�Ed��7�����=o u��o�`��/�W�R#սsx��"@��c��Y�J��=�+�qȡAk�3�.�*5enӅ�;�wnI�$�.=@)F������/+�]��P��Oc����6�m��[���&iKo�,����e͐��~.�ÞKu��PѺ��7@�f��g'zA������E	�������C N����v�u��G�ڹ-\h�����A׺��x��j3١a>R���)���-���g1�����+���F�vͿuP�V�k���k�< m3��ܒ-D¾�L����k=����������z�[\U�<T�))��ч��c_v�F�U��mN�4ܛ���/�W��%T�oz�����)1���-n`��PR��t&	��+]�PhqT��_Ej�/p]"������!v�=����iW���&g%jx����<���nE	��$�. �SČ�n�<4�>u�
S;�[>hY������8]��ڴ�(�\)�������:uD�,��栬�5H��2��2�����r�߿L�v����^��iJ"sm��X�!��1����"����v%�d����&�4�-�(�S/?��Έ�k�~�h7;wo����p[���mCQq�㚀Va�\)'B�6Ė�@[|9^�U���f���=�>�d0��h٤m����jT�ߐ���7�E1Dqv`Nb 1�]�s'�Q����1\:��dk	�|[����d>X��xȤ���0���T5+.�r�1����~�����.X�+�(�&�'|����F�)Y�3�}lW��ꕯ���\t=Tb���~لȤ�&i��j�Xw5��#w	 
ں=�m�����g)�[>o냑�gIw��f��*'W�p�� �
���\8�ս�X'���g����e\������(�m�����5 �'٬���\���n��9d����h9���p�쮽�ƨy9�B_��N?��a�$4�@�~��\VYU��K�P�)�Y���� ��^���u�:H��+�29e5[�j(�����0������m&���d���t���V �8b�N��whe����g��G�J̲-�}��{v[T�*�� ��mm�ۙ
ǯ���G��uy�b�a��]޵�4| yD���W��t��nrȓ�vG���E9�1PģtR�O� Lr*�d�o܄�Nd�Q��"l��a�>���'6{�zoj+:U�-����S� �P +�]k]4�(_�L�b@6�W�t���1�#���Gg����82�5
����VãbG[-�= �w~���Mfi����	M��B.<�u�_dz����]`?�}���L��GᅥX��6L�4S�k�B���Q���{���4��]_.�iףV�2)yec~�e �m�3D.�Ԯ2��VS�o��^3*��w���,0Ȥ�Fe�)���u g������`�,.��P�?�ج���k��Fc��,XQ�mdM������B/�A�G132�!�p����F�\�8�������>�)������8�T	nU؍��>��K�����yM2R��A���5����� ��p$��@NteH���n�[�4)d�"���0�[ǀ�Fw�E���$+�Aȁv�p"���MPJ��8u9�vYb��$B�_ �Q�`82Tx^�a��lR?d�Vee�胵&���J��J����fj�S�}q�P�g�Nş���1S���9�m�����=e����NZ��?��� e���y̡])�}�d�g;�E����6�^��_�<� �,ᇫ������ԟ6�O��9���"��C3��Fk�Æ�k�2!�A���v�g��3)�m.K��x��Ȝ����7��+c7!���х�l�Q�p����$�X��66�
�n��\p�0��8o�~����[MÞB���ܛ3��G1+��F�d���?.؆.��v��@O�4r�A,����p�>��.�/a�cɰy��cAs��N���߃����r>�9��������6	uI�ت����T��B����7 �/%z�X���W	mٛ�`�?��b��Dt���naS�y�#�ߏ��L��Z��v�c�)$ ��粒������������Wf�;�	��k�/&��WJ�MNsJ�*�����O�}
�0�!�
�ԁ�LGE��C~"O�5��P�lވ�:�tB4�x&Aё9|���)�𹢩Oq��n0Y�+�b�Uʊ���%b�W[�nɮ�f��{�:
4i1���EE�nh�U,I�����w��&�X��sD����;<9,6p+_8M��-"1����Ϩ��xHp��lO%�C��b�c+�	Fͤ
�n�`lc#�tMx�M�d �u4ń��'!����'p������V�9& ZQ���90@2�pK5ٓ�'�:ݗ� c�v�������%\���ܠ��'��#�b�Pb_�Q�a�S�#�ެSOs>J�eqd���/	�l���¦�����k(��	����9g`R�_��ܣp���G��ڹ9�݈�B�I{&�L�3�!A�Y�)�nu�$��+�aY�x'���O��ڵ
9||�ǯy��>}A8���o����:H��֏�4����pn�+ͤ�sŀ�r��ήz�V� �0��	��ni�g��"�IX���$7���~lZ�J���!p`�tD\�H�bDuOJ�H�Ų�1�њN�����~୏�/7�MY	 �B���Ly9�2lH��[��ӭߒ�Ұ!l#����W�u��$�C]�;��_y�o6�|\"��~w�~�n�8��QE$T%A��ȭھ4?��1���Ѯ�vX��-���1'��B�搅��q�a�{r5�E��	'��ۊ���g�AV+�+3v9�&����JӚ �V,ٸ��]��������ƨ3p�D�ڒW��M��Ϋ�ecR��r�\���|ǽ��5З��>��D���{Β*���S2B�����B��@�~mm
J3����E����)�b*��5���TKyc��G�ޣ?���K��P�$���7��ٮ~�J{��������$�2�T�XTv:(�ss�=`��ʲ�m����M�u}^�aRS1A�:%�蹮�x��=܁�)-H�''-�\Trב���z�/d��M�$( 4�h�8r�qv ���LsR0�K�D�ѵgٿ���ơ���f�v��sa��p��8B	�`�=��_�#�B"��C�[��+h�/kӊZJp[���	��y�nta�o��G_�5ai�N�u*o'ڑe����ݎ��7���M��-���;K�ܐw���4��*p܌͏Ɛ�衾���,��4CP2��9B)rC��r��I�� L�Fvͧ�v]�����lH9	.�.�r�>��A�+.W������^L/� A�\LW@�s�{=6ӑ��I1)��K"��7�~2����V
��<4�7ku�����T�c�V��s7N��e�8W�?�}EB�Y2pn��RQ�5I�פ��<���3�t�ݽ0d�Qy�͜g�5�PUz�Z�	��u "�Y��������t���!�@\�ঽ4��LEU�<8����/�K�$��:�3:{��a�����9`�����!�" @K_o_z�?Bpu_?�XDG��ѷc���eh~[Y�,� �_��4�pA�[��Zq�C9����P*U	���=�W�����)�|��Lw�&�F�˵��z�3�./	·�2��C�V����bD4��Dԩ��6��U
MCqao�c��s��B����٨���ҿB��4SL59�0�׻�����^#����fR��L�³�������OT�F��8��ɊǷ�y5W.�8õ`wɵ� ��xלC��IQ�MVMNxP	�$t�Ć�Y}{RNe0p���`��5ӷB���� �I�
��wD�}���lr��G	����}øf+��qн��r���m�&K�JK܍�$�n6 �rI��t�y����a���x�u2)q� ��B�/_g�s"i�"�R����d��`U���@��CK.�-�wW,�m�������0�s6x����ȩ�z��Z$���{�q��8��5zN�m��}�<R*0F�]i3Zَ4OJ����]i%��ɕ_�6�g�?��5�Ë2"�|M7��uˠ�!ढ'��� ���9dk��y�8��C0��)�WB���n��q�����/��+���WCbP�k��L4�Ml��V م՟�\\{�4�d�0���X$�ԎG�e���r�)����W�v���?��X��	s��b�� ��
,�J-+��-����Xn�볲ͅ��~����ܴD01ス9�ؐ>�
�i�zl
֏�N.w�<I��'�
�w��so�ͯ�Ը��޷�;J�C7�1h��������Ԫ!�{ZXr�y<s�\*�{�����~X'�l%��_��]�f�F]P3�d�󟚷��qtG���*��7�'2�Ok2���2�����i)����Z� q���8s'�é	z8���ȼ�­T&������ ��b/@�C?#���+u�e�9���n+�����8���KV�/���/d���5v��⧉׳랹f����Ϸ�U��6��ĭ8�)f C��\�V��A䵢/��$�o����Be�wo��Z;JٴJ��g�m���<ޘ�:����g���D���&�����yj�^�x�>�#�dLZ�\x]�$�r� g�V8Iu�f#�c���pY���FƊ��e�;��k����q.;�]_܌�杹D�D`�o)c��u��z��?k�j)(�������lg	S�R�nq�ҮMkg-�����2�HM�:yfB�p��K����h�gS@��M�~��L4@� Q�6x�|�H���U���YW�2��}�蜽���ݶ��	��#��f��9��[���!��������7I�ޥ�@�D�T��%��.ONn��O$_��PM��u��K�'Y�u�0���QΪ��$�`�Z�\sܵ5�8b�.ҔwK�av'�����~N��c_�?FO�(4@��׏RVm�P�/7�s�1��L��%s0h�!�y��+��wo���2QC_�X<ԯ��VUM�#�%�]?��Ĺ|�D,�ͺ<�����U,<^4�Nҙԏ<,&v�z�uq�|��Õ&n�_��+C���F@z´&�)ڴB߅��O����2�'"��Ŏ��1A��5r%�q�RɊ�0��kQY�I�Z�L��' x����KlᩡؓZ�!"Ӹ�V��*�L�w�js��U���7q��زc�y�`������a��]@@d��tDO���,ΝiOKl�����y�r5�e�LД�$�V�ȋ�KV+�m-�B}�������D�;]�!o���Pء�F)1���d�\g�v�R�Ga�I%��R�����N�Z�O�i��W]������:i�	��q�i�t0��0_���R�����5J0¼ql�E1�Ӭ̊V*O.l؛��_��a��X֜�� R�-���feZ?�+�-�����dk�3]|X�F,J"A�S�֮ڜ��=����(m�s�m�,����c��.���ԛ�#��V�-�o��\�K�~~E�W�^yB�|Ϛ���|
 san�r���Ѹۋ�7{$U���P��͇P����������ӄm�[yO����J&��T�gd����)*�^�*�W}� |$�!TmQ�e�c(���MJ�=�G�.��<o'?��{��;����>��Xo �¬0:EA�t��Y|笈	�p�g�To�s��ie���ueF�Pq�c�(e�X�*6��z"��ʇ^0�^5�� �C=�I�Ama�$����8�I��>���Ռy�+��m�(�Ckވ(�Gό�E�W�@uqq� ����o-�4Ble�k��%�7xNӜ��W?j�3,Pުx����[�Wa1?y�u&�C��m��7�e1�[�<ύ����Ļ���UW��!���N2Q��t��q<��&��O��>jj�y���4����A|]f�Z�x�f�rH�!�J@<C�r�RP
e��+�a�)D�(�G��������CT��{�Td�m�o�uMfqۤH���&�j�;k�
�>O���hL?�������ߞZ��)����=Iұ���N�|�ivƕ�������X�Ӵ�T	�/�7��B2�ƿ���-���B
���=y�"K	�T��~ăR �\C������R(������H�.�������o���O���lzI�Jd��>w|@�q`�}�U���t�iK��������n'��4��\���0v$�Op�]=S^v�@��4���� C�a�vi6�MN���r9 [Iu������������B�ձ<��V��+�W�H�s��w� �Ʒ�B�c"�;J�#%Xp�įHy&q�PGy�cC`CAz��41�g2>�����i�0H���م�,��^gfX��A9�M�`~=l�2.�?�*����ۮ���ʡP��u��(uj,�	1�ӈ���U�ݥWO�<:�m��@���WgP�/�fd��w�bx�c��1|�(����d�O�U��(u�(�e}���o�iY�'ʈ��`J�$�)1N ����g��S�,��ވڤ��'�Ȥi�eԡHҳ�v�9��.������Pv�-�`QZ�+y��q�$L"�X4��+�����C�?z�%}�"'�~R$�ȱe=�H̘*N利���7���##�}L��=��xb�ؠT��L�����(��M���ԍ��:���K1DZ��E�-g��1�tcl^���F���H��ٶ!�*Q�2��y��i��A�8�ͮ_U��{N��+�4��'5���w.I�$�D0c�`������-�^�4,@'��
0I�&
g���'�Q��rzS�>a��E{�(��Ε�6��r̷R��2�-0`("�~Џ��8��i���HI�Q _j���ǡ��<T�噢~��3��� =�H �'�p7*���!������߶��t�����'_a��yM:��v`���@XIs'������FQfR�.���☕[�iՇH�֛!4��J��(��)�>�z��d�K6��9SB�;4xG��%��A�$�}����U���h'�H͋iX��z�*:�9_w�p�=�x���e\k���MZL��� �K�*J�~l�@l�1N��� ֏��Pq�P�Y;U��P��'�:����{B���Ae�/�d��@I�|"���
�%��!,B���<o?�+�H"y��S�7'b�/ļ0��^��t������d������2� �:��3aA�q�٥( r�2(��^��V��_��#��h:��ti^�}�>�4�y�l�t�b[h��ĥ��\�)�G�ĥ!
���u��	�[n��ǆb���-���6���Jy媾�訊�)��8�����_��ehҷ���}����\_+IZ���"�u�57ɲ�d��c,�LjqtZY�\�-5�-t� �e_LB����xr�Z��*\�L�u���϶��S���J7����p�y�-τ��`%?�L��U��L�Geb\�e7HsPS�a5��$����R���p2��ͯ�M�w��{.?a��q�}l|��(y�����j'xIl�%p���(�<J�v��N���F�cAk['���W������v5&p6��i�c��,(�IN-�2�Lo��N�6;��4����Wa�F:ς�n���g�|�G皣%Q�G��^�~�������;��v���Bv4@k�!%v�b8}T�����уH�,��	/���ޮ�ml�5�s�y��^琽�e�uq�5�S�Gl=#��@�ӡ��]���x<[�����g��hi4|^�R0�L����96������r,�C��.5Dtܿ��I��n>Vp��N)�]���l��s�.�q}�KFtcF�M�L9�*�A�a�z�;p���<�zrK�
�
lb��$,<�(�O=Q�t�O I�0馂L�C۾�
��L.}"��#!z�H$�
�i�lgh/���1�<	 �q�ٰRDd1t�'f�6�7��K�ނef��V�L}�y���J��4a�_>�1T|r���\%G�x�-ǻ�eg��ߡ�aI0��mD�T�q����]�B��r#Q�� ���`�q}�}��C���g.P3��,�M߀�$zcΐ����?ʮ������ʚ_�������]@S�GtMÑ#p�@[����z�M�׼LKӜ��.QѤ8y,��Tg��0�kZi���<��.��Y��_W$%�o'7��GGA/c��+Pp֜�"T���d�6=����b��Vb�bgB��G0�_��^��S��㼐w�����s9���VH5��q+���ˬ����z�'�p��D@�M��ս�±�
`�0-��Q7v�޵�V��ٛ~� %Aw�8_>�?��GB��w�R�QYhP��|2�����]��&h[:v)�"�s��<C>CW�87�:)��f�&1���v�Ā*�I�������\�#�PaUZ�S�OW(l���˷N?1滯$�G���q�4��2ODv��D8�h0v;��8���s��Ƹ��$�:�\�S�P���^-4��f��9����n�Ƚ���v �^h�X��[���o3�寏�x������%��+HB¾��z���{� M
gq��ř��%��_\�-���՘7�Z�����!e|�m8ą�h띵O�d�_�^ L\��!�T*ê��wd� ���m{��F��GĲ��%�E���"�2A�8���V��aƨmҳ�dJYV��qu�������=W�V�f�� G�=1�w���@��r�y�F��ಗg�`ť5��+�����=gߖ>�}I��#_��3Y4t�'eJ+����cv�d�G���(#���2���R�Zp��Ȳ�͐�Ѭ<��18��S��x����C_�6,,ϥD��!��H�!��9[$
���4�Grj�)��W��p��^����֢��0�J)���~D�aկ�����I��:�K�ČG�Ggadk$�֧J�G$�[��y'd��*��)�5"����n�����Y�6��h�Jd ��=t���j�����B?���~����8�,���]���o8�o�Q�1knN< IM��?�N��w�X����`�@����i��0h�)z�8�~�@��~���h�5�Q6�#`�D��J� 2���P�b��C �r	������y2쫞�'�� �x�i�\�tYwd�0.a�T�����ک���q4(�^�^0W�:��<��:/�HF��Q�mν:I@��_a~��R�uc���Ӵ�"5��WQQ�KP�� ��Via3�)L�j@�Q��i�N��5Y�8��Ι��.V"�n.�8����kܶrU`
�a$A�o�����UKzeL,��@P�R�[���,a����a75�����eき{đ���L-����q��ߕ���m�}��G��N�D���̶!F\��6R{�OA���|�&�ʑYLŹaN:�0���sE�؋m�`'���4�h�Tv!��7?��F�ŉ�7Ɋe籦�������{�=�/9J��1*w�-8|�@@Lv�{�W�����ٜ�b,3���ɷ}A{nV�T��2��d�F�x�Vu탐�J Jf�Ekw��`�9�i �^A�QִJ&��� ���n�}���Q
�Iu�&!BF�q���g��X�9�O|So*�6Շ҅iB�!��Hn���K?aU�[K�/��� C��*���.�aZ�䄅#sfK����x:������9p�̇8P��~�9����nV�H��Y�>����qGW�)�|���e48�5�C�py�B�bnٜ9u���Ն�z��)������� �s��΢{�Z�Q*�� ��Z���QK?����S����Xƻ��#.|}T�~x��9�b_V����jл�L�vL@>��D�ɕ@��~�5��=e[�|D��0���kj�s��֓+�M�>R>Jc}����w����m�G��i�+�1#C2��;�Nw�[r �C�[�e_f)�-��m#��	0}�~x���z����*�R�"K�q�m��njLJm.F�C��ȑ�{{��2�q��W������;�K��<)�C+�2���v5T��N�Ja�2L���5�u�}QN�����{#�=e��{��?��a@���W�0��������/�
�Oq�䶛�,���Ue��m1Ǵ� �X�+O�r0;��=�H��=�L��)���+�޺�1����T7�J`�V�/��q�b���lSU�E����3�M]<'�Qܦ3I���,Լv��i5���MifZ��'M����=Ӱ*�^o��W-�Lh�.J�޾�����Tr�H���B�jt��dq>X8|I^�p�Ҵ�]�+�<��7�F�L�w���-��|"	4݉��ѿqJ_��2s�:8	�����ە�m�ͤj�#l�G��R?U\���������4���c!��S�έ+�{�xr�X�:��}23Rt��<6z�r������Y�#�aP�7���N��
c�, 
X�ܦ���
Ӊ�v�U5��� ���-ٜ{�@�A�3!<�ɰOc�
�9��P��G����B8N�.I����x������_��k����8��M`� CZucMO�	����^���s�ׇ����^�i��qgge��	���/mj7H�g$�{��w����Q�'�ס�?�-/�9���e��U2<���B��G+�#ߚlH�n�Կ� ��JXw�������I��,%.�������#�"�����/���>�<�h(r:z�p\N������}9,+(N��h6��"��fn�lɽ0�[
��#`���<`�Pyí�Q�ƹ 5�i\���U�����o ��Ћ�ȭKԕ�J�Qa���S�3<�d�ԯ����Z�ء�g�*7Ԙ��;�M|O���yi�����2�f]��o��:q'�"`�[X,�O@T-���wpW�
�J��q.ēw��5a�c���x�.y$Cl�"YR�%>B(`��Y�Z��E�0�{�B�4�k����g+���C��jR��_>�S�9��Q�Z^[o�7Ȋs
R��4���Zd@���=��$�!���)�ȟ��9LV;Z���͌b=ChRʿ,.��~����+tց�*���%�F{y8R�=WN��M⾁\�kɃ�w9�\�Mm���1�������Tcb�{%Ѹ3�uq�'`����ʬ��u��L�ԅAE��"��lW��L��|Ų�����A~�@�X��ݶ����@X�� �a��.>(u+��[��?#ΑT�����!Ϥ�B-�B&(D�V5�7��gř����"�����-�B��
��v���&j��n��+�c�ɦ=v����!���t	+5 ����+Eq�븎!�Y�>��؝ 7���sV�'����Ul8�M�6+��s_+�r蟞��-w=�l�D�>��vM����a�A���E��Ȼ<¸��
��"A,�m)4���{\�6��|i�A�Fw�q=*s�6�2���)ѓ@����4���UQ8�a�i�\���8�a�x�/kM�"I{:����Xy�񋽓�x��g������]����n_j��/�5B��uE���g3�0�-�_��f��I0��C�'I���R��)H���z� x
@Z��n�,����J�ͲX[]!�H�L\�a�b�/��P�WϜ�R��0�G�YP�����M�����퓰�7�}��ͭ��&g�F7��ޮ%��)�*�C눜,b��K��7���K��.��c�������@5b��(�E�`��@=�nm�H�&����"՗^��b�Η���]�kz�6��0�v��%�ir���HE�6��h`��A?*��9��RcT֬)���yF�
�fr�*��3��Ⱥx����w������\}�ke��W�'����=$K+K1(�b�vH�3ie�۫�Ir ���CSK�V�P��\H˫�4��7���*i��"w�Q!#M�	��T[)�&��a1kB]�]��y!]j̚��0B]f#�i�F�Wǹ@t�I.� ZҔ��䪈��X(q(	+o#�	�ff�����7��v�f���'Y	o���9'�B��2���c�j���3�;��|�}v:�g�tH>���L�U�a��$�,�a�AV��������mH�4�����-�������cku%
p���#~g���l��B�8å�3��K��+�|��-��5�2��a�R~>�:�hy�}S��<z.*e��;�k��PP��Z�(c�A�424&z<R	�`]y��!��,�Zi�w����2�w��\�5�=���?K\���9c);���T�N��Y����a�R���=W��+ݒ~�,\� WxRq ��ί����N���7��}��,G<7�K4\=��
��nZP]~6^�q��[i�{vt(����%
����~Sq:;�ēv�뱂�Xi��Su�;/)��EL[8�+�_X����2���������9�r��J�)c��pn����\��E��<��n�M�Pm�]ϒ�/�"EX��Vd���;F1����d�R g�2P��4��G ��P��돠��A,eYͷ��&�+3U"�V
��2���j�'a$ܞr�B(&Z���� ˶��Q�oq�@YX�W7�6G�t-���6n��:!��6�go,�,��\��k����sd������M�,��x�[�(�Q��`Ս��nQ+����>��(��nh>�a����_�Z����"�G?T��.A���Gt�|�r6H��f��*҅�Q�ZgA������E�l��^����h�ԈZ�WX��ò�8��CW�Xh�iqȤU�����N�	Һ(w|#�K�s٠�[�=zpԒ���D�N�~h�������S��i��$�X|�r:��>�	�U��u�%4�ZS�a!k:C�'���q��G�J��;��x�
c�L�w[��M�kI��g��
��d�y]NA�bȩ�v�׸b��1��y8ۚǱ�M�YKj;�sw��� I�ÈۈU��ۭtW�Yp�4��1�YF�в�Ӌ�y�Ss����)�D�j֊D����.�x�v/��E}[���I�I��U����c�!1��ܲ�[F�wt�� K䊷��m�G�|qH�����w�]Ω:{$+m3Ǧ}ؚ蠊�MW<�-�>b�;Hk�"e���3��W��R��	��w�!�?9z�yR��R-/�J�3��z�i @��`�2j�����b��R�Ȉ�9�h��Ul��B�dp��b���2(#\-�o�k��N��[�����U�VH�94:{��<p��Z&�:��|Յ�4�ޫv9f�|<Q �ެD�\hR�9��+ǅZ��\�fn��0Ui�=������(bD�i��	M@���_��k�vahK��/	��DقA���֚H8O��N��-����
�NQ3�n��B��g�Z��@k�oB�0�V����H�bB�^�?$����VF�.h����'�]`��S>]wB�$���5��j���))۔^"=�O����Po���7ma+��ن�|y�~�� �F��7���E��cMˣ��۹��D+��`�k���N�K	���bDc@��Ӏ�W�g�y�Nޒ+�|��"��z�i�E��F���?�=vvB���r����a�P�}��t����>"��4���8p' ����j����5D�5�L�����9�	�&{�?�r�MS�	L�O�B�H�)5L�xB'%������7?����X rM�����:)��.�n<����2��K��勳�c�`���X�z���_�g��q+��!�\��|t�?������"2�x`Ѽ��[�Z���|��cy~o�&Ƹ�����#��ɩ�КhL�I�Wk�󍕘e�'v�b$���{�?�+-�ȩ���,����ަ�]�����룚uqk��Y_��u`5e����*˼m��0^��4��b@ܲ�w�$���<���";h��aL���N]"��
�@�`?L�����!|��NCn;�C�P��W&YD�{H�FdV�:�ap�d�s�8���b�����+�~S���Hz��&E��i��ي�we׿	�$3j�滐�f�	��PG��L{5Ԟ>�xђ��} oU��˃�ϣ%F�"�l)��/F��o��`|�N?�����C��V��녔N�y����z��1&���C�̘Q�\� �ҫ��H�q��x�����jY����:�貦�o>ۇ~�3�Z�ш�G�%����*LI'?a2O筒Q��O�y�@�+K���S�&�GsVn�~&��)A�Y������1���Ԏ
��^٪v�'�o8is,���Y�0I���*�\l4���dZ��u�GK�c�8]R8ǘ��B���k�����;�<%�.5_n�E-��<�(��F����>͚L��ტNX	���utQ��\UD8��kbVѵ��^�e�~l�|x������HU�:>F����k��9�L�2]'?\9ė�_fq�$� �V�p���UV�p?�[5ef��[Mi./�7Dl�PW0�Wp�<�O��Q]y�Y�i��z7P�+��-%/���8��~�ݯT�X:uͰץ�l�F�X�����l5M�$��D�	@��x[�`��8�$�u�]�u��,�N��̀FD�()����\�WG�)$�Ǧ��1�#Ʃ���^�qW��d<'����O���f[�i;���>7v̴��i��	�/���w�t����v��� oޜ� ��F���j����]~[i����AH�Y��4��eE�q����H!�%���4�#��Eh��J7���SMY�p���x��/���8�|��h�ܯ6�V��3	��a;h���OW$�$-��4nO�Q�B5GeK�8�3�U.�S*F�7 sD��Q��zO�����B΍��q�^EO�����V�/���� ��iǒ|�� g/�A�}�F9u'��W�Y��@���D��69�&`H�b��$xl&�m�(�˦�C�)��Y�0�H(�_����;��#/���.�yK�Fv�6�
l�9�Z�'$�А���"=�U�����.Y��j�|��Lz�������h���A6�x^nu�a^�׉+��f�|��C|ڇ�-�
�~|�ˈ���7 �7IV\,~T={�h���.*�]^���Xyw�۠͜�`>�C�3R��%�&;�hE��Hi����B�A���ވ�j���+)I3��=S�z,�����M�$w�4�'�k�z�A�Du�?7X��ĿԽ�F���$XMN��"��^���b��h�(��j7~��{�Iwf��V�����������{�6R��3釅��UV
�V,��1@�Ů+�̴ zP��4ޛ;L��O�9�`M��"S����3�����ܩgl&9��	��,�v�bb�k�h_X_��֍�ӟ��n�_0Q9���w���i���kfI����0�����`�
�=��'N9j)G���c�t'0�JA�H��0�X����	 �}j8��19�"Yv����;7`j���DE;��X��eS�`}��+�I�Gn��G����6U����Ď�ڔ�?u���O0�-P�  )��g�È��꤫F�Bʁ[��sQv��R���ܩr�u�������w4�#Pؖ:5��j��r�
��ի�vw����]�D��)eG��W�<gr�A�5Cy�'ż�ݭ����DjKd����M�V��n9).7��i�����6��Id�S亏/w�=ʒ��/��+�FD/|�q�#2�܌�-��K��7����䍍���F����2����C�C�V���of�6���Mg��GX�&�j���&ĘX�Y�)�K� LsM�)��{}i��7��C����e�������M��JG�=�?�����4b"�:�DI�yt��;��.;U�M�s�Q�ت�C���X�B�\fc���ԯWs\�n?Xe�&	�l�&����SaF��D .�س�������YM�	���}SGK\"�����_?e$[�-[-OP�S���s���c��9��kT�R�yL����
�ɲ�!�e<QZ^�c�Ce�!����m�fy���N�T�B��=��]:�b3L�����u��i�Hzx>@M���񼷿_�������`�0��ID)&��?�HB+��"�j�$.���1�۔ڌp�+՗fgQD�:+}���gCI�FDk���\�U��>��1�o�����|����a8X:-zy��^K°�[..�ͧ�A|�����t���8��5)��7��4r)���Ġ�TY,��Kn�/�ZL�<d/8$KQF߱���Z>��[숚�x�l�ǖ��Z�M��8<�2'w�G�O�b�/��gn$��f�J7E�)�C�M���z�ޤ�[nws���cfϗ���eֱQ�����D�+~�7�m������4E%��3�g^J�aA�/0��#7Sz����>S��/�v7�����N�����w��vY�W�b9O�%�3�2�!��_������H?�&zn7�f�1WG(8��B�M����{�@��M�_���>�s�:V��8\n�Ğ����V"�VUz��C��O�}��q�� �t~ˍn&��l�f�;�
F""�ŭ�Xb.�-O��y�xo��p�<��ۿ|��T��IoL�飌G�f�T�����v���=��)�����U�ޝ��(��$�K�VD7Q�ɱ#*n_�>���I�cҷWӊX�,���D݇�&%�����
�[���a(8޳��^�+��l�~V͘$�	 :�
�JҶ�WE�,�UW��${�k �d�!Rt�x���o��+�DV�n�X�E��0K��w����0��� ����Qj�g��vg C�O��r&�ig+����͜�a�$�Ĕu�(���;���Z�S@��s��	 ���\ ��J+�pz����i�-������m�ΘTb�-���X/ JRf8G,����][ �$a+�W�'aq��`E�u|�ld�Z� �����m9���iW�ݖ"Pw>�J�q��QS�`�d*dӧm�(y�K�#�v�D=�=��<�\��X;�-&B'��!X˴gVq	�c��ҫ�e����}"��/�z�f;8�.��c��L�S�ۣU~=>���}i��~�}�_]�ٮ�9ǿ�
Ȓi#H9e�W��cF$�_�	X�<mN��`/:+��#�ԥ7��a�M�����'��+�0r,f =k�,W�p�^�F�p�����7�-����>�~�H��ɚ�hx�ޡ�D,QH#"w���p� ='��Njn�\�=hH�77�э�Q�����!��j�U~e��<�5P�X����nV��'r���_����9�伢�Y���0�l'ic�fN5M� �R/v���Cʇ�*�U��Ѯ�+B�쩁�]�(�~�g~z-{\ϳ���a5{0���)�n)�r�n���/�QJ��Yi1�Wv� ���D�D
����4���U+#��S��S4%c�ޅR�v	�̈́լ�� 3
i�D�o���*� 4�~m(���A:o��e�X�݂^� S�v��6n�`�NZOΞ�ҕ�*�ۦ0hkqU�J'X4\�h]��_��Mbၣʍ�M��yK�V1�9�F����T�^P%$%!t�dW��R���k֔l�����s���c��H}{�Q�"F�+�f/D���z�<SM6�C�%����B;��'��� \,̉Sxۗ��y(i��L1�l��ҟ'� #q"��_�A0�\EU���l��b��$�ʴ[�]̕K� K��T"{Y^��{
���a�Ȃ�Z���\~BF
*�D�:��S��0��oR)�O�j����ZA��u�P��['�
?�r����^.gJ�11���s���T��� �ifa���8����~i������~�4��B���� K�.g�c�݁�$��V�2Y���Ś�!P��um�q�09��ă�tV���J{}Հ[8��g����u��z&���;,�lOxjA�BOt��'~.�)-4$F��4�t����UE��/&�tB }��&�V�jqo�����r����^�
sʑ�K�V����A[����ä����K�����T\�_��Z���#�5��v��G���R�C(�}�A��h�a%w�}�t9Dy[��4tM��3���e���p�:S���h�~�"����
&�}�1yv���_&=�)��j��g�y��輻�m�Q#��A�~��]�"�m�%πI�fB�y�9�%:�2<�o�B$N�����6�q������N����2�'�k�9�Pݴ�~�(����������@/_��)�z��H!���ie��������ͻM��u����D�*�+�30B�$��[�UQV~��f����N`�����	��1�pě�Hw�W mA���%�+�&C�X�X��e���&������%w���H���z�_������\�>H]"��!�.�Q�������Т<V�w&���V"���o5��\��@��4 (D�>|y�-}5�!��P<U f8 ,�d:��c��D�S�:Q��N(w�3�AM�x[E��a4ߌJ�����W����G�*�uEj<<��Q8���J
P���N��8%IKQ�3�����^�mt�i�� `���p8�o�2�v�2`9�����^����y4�0���$tYq�cK����>��58@�Gs�T�-4���(Ƴ��^�G2􅭖�'��}ʙr�m	�`��I�ĉ���Haր��>�zJ�ڡ��o�PÄ6M���a0qg@��鮠�pԭp��F�}1�R5a�^���	'Fzy� ��iM�P��;Iɿ,�y��l.D��S��&�"��&��S��isL=�8�����E�L�D���u�	&g�ɻr���
�¡5L�Mjb���.4�J�^�6ݧێ��-~�0 �芪�G}-�l������9�\s��!i8ԍ��UeQ�A���R�I��9�y���+�U��2n���~���#��1��1��sQ��ze6E-|j�g&=��Q�Ϧ!`�_f&���gu�W;~`4΀!�l��}��	}v�pV�V�c�C��JqG���&VGОwr�M-9�)7�!�R,�J�J�����3��k��sQ�z����u�1�Y?��@��X��9�3{��xfm�ߝ=�.W���[9C�Px��aʠ>:�fܵ��
���I��c/|�λ1�Q���O+�̍X�"����$��pM`2ŐQ^�<䋘�.��T����Tin񹿯~���1<��١*e�$�%QxG�L�?{@�%�'9���[I��<�d�mɴ�{��7y����%����3I����聱�YC�x�J�]����C66�1b��e16;��m���q�l��gF���w0�N�%\@��bV��<��B�\��I!����(7I�W0��&�C=��l{��Ĕ�(r�#��I�%�P|�w��d�"��aL��N}�1��4t�b��Sg��/�s�)l�"7��3 �P0ͧ��6�tԧ�=�����b_{R�e�{�J�ڝ6�t�cT����׿�IOTe�v%�h�cEE�^�=���ǿ�(~J`��es��n�P�83"	��B�'5��n�E�@���"�E�XG��#(��EU�g��ӝ5$�N|��O>�pD�8�ө���A�_2R�(8�j&�s�^�Q^	2��C�K��ﷂw��R)˺�	��'������e����F��/��S�/�@	d˟�˳"����>a��I�>+�Coo�)x�G�Hg4�N(`�~�O�R���p?8�������G]���\'�f���]�H
t>�Q_+h>I�0Pk1j�j	�OZ�h͟�HK��Z4^W��jFh�~m�4�|�;���	AAi���Ro:+Ǵϔ�	z�����&�m��g���%�fd�d�ëZ�دH�I�&���ٯsa���ʲ`�58ڱ��=�4�hmt&������h��X�&I2��^��G��g���˙)��ə�ͮ�WuWO���Ӄe�`Gu�yʣY!~[�Gr����Gs�.!	� �N{%컄����P��[����k�Z���z��I�/�l������{j��u6��}�� ݹ}��/��}��e*]F�89�Q�݀�	-/>�eqφZ����;���p��g�r����6�V,du��幇Ǡ��rL�����_� � .D�o��tT�MC�![������P�X{�O��a�����{�	0��gZCP�JƆ)q6T��#�}��y�k`7��#rҝc�������U�b)�C���{Qʡ���Z��C������n�0��1�g�0Cf��s��^����7?T:=�����[�[�����.n37�ȧ�Ά=VO=m��A?A3�3�2Vכ&��W���H� /fb�3j�#3ħ�kW�������h�fL��KC���3݀��ԿFCw��ŉ����*>֨F�Ӌ��A�m�˧� ���� d�恙8D����f�
�&uF�mN�"�u�|Z:�;���A����5��;Y�Z��& ��>�<a�5��1�YB��l�V��iGD3S�`�����_����i��U+[p�'����b����ҩ0����y�Y�31��O �&#ft���/�����F��4n6��Oѷ�C_�ܿ2_�P�.+�<���#�U�==,��bXh6n��%rH���?�-���8~i�q��:B{^�u�pDx�9]�2H�.��]���9�q��ߌy/@�52�����'��2�E�����?�xA@T%��!��~�/�L2�Z�_��8�x�S�|�p��*�{sC;��ӭ�P�E�hK�}k��Ä�ޫ?k鸫%���c��9!hgJ�c��ې������Xw�f���Q��ڿ9Cd1�J���Y�$�+CNˮ��O��Ð���"�MpʁU��猩� _���.JU0{��C���ЕO�aX)A5��e�Ip��Ў�`�*+�B�]�G
W�`By7	��q���N�ų�-�dn`uOrYE*��.�vb�a.�D9o���zʙ��OP��{w#��F.�D��su�L�w.�i�Q��Y1�JWIdS�&ӊ.��u����3��ۗ�c�B��S9�R-R�9퀪��Ί�]�4��վP[��ˣQG��fS����^:
j�W�P?�]�7.y�$v��I.S�`ԩ�����]�H�����-����z��ф�C�N�34�	�ӈ�ko�üV���D�}L��D��n����j]�&|�v}S:���-���n��4��f��M~��i���T�-�>��5�`��0�8�=��	h��̗n���L�{�dY��`�Ll�!l���^\�J�<Y�����v�H��\�T���M��wa=وu���$ >�0����]cq����zE5���|e��,�h�h������O��r{��륱��v�@*���)�w�
�91��,�kP��_M&�_rX�g���~?U��,���Z���5]�g�vTw��,cWڝ�HY�o����a$�� dͣgC�n~�n��������-G�1���\n��g��]�*
�c*V���`k�������Ĕ�>�]"����n^�N5��p��.���Q��"�]*�c�UУI�%�'�.?��3¡���&"h}�F�Q��E����D�����=Mv|�7����n� /rO���w,cقObu��)���!!��J��D�%xPm���lXrL@n�F����-s���hD��*���Yz�Ķ+��v-2��rѽr������M�,��Nb��Oe��vk��q1����PAzm�\U�� ���!px���6��ƅ*+p~�}!��I@����A��g�
�2�۸؃�[�K�$SL��?�Y8��)�b]v�I[��n�������_���{�$��*���-|Mݴ��-K
9\&8��T�(�n�̥k��̯{�'�Z��'ۓ���qs!<��9r  ��5JXi�>w�Le�ý�)4{�jL����m�3���a5���a����h���)�=�2�i���_����6S`���R\T�,É惰þ�ip�;$(2��wsF|���=�"�zȢ^'/1���r�^"�r-��Mf����7:�@	lE�'�*�l*#^�<N�uk@�\�u��E0���b*�0�ז+ZQWP���m@��0~�$�����r�_�`fvS窹��$�Ԟ����l�t@�<ǿqHg#}p+ͳQ��c�b5��J~��yiqx���&���\d8�"�%{��n�����r�-��m�C��O>}$�8�����	yl�j<a�J� �SLԭ��稜��Y��jI�M�v�6�𫎂����[�m�a��0�q�ϢFs���.�<̥������cq�Î}���aD�w)�WQl��\�Ә�3��}e�9��i�1��s�	�����#���:�t'�AvoC�	rh�//��&����q�y��^�M��&Ԥ�]T�e��
�Am�P�����}��Zy������Q;bC�����&��<˳\�� �s�{�i�����Z�{�/�f�UQ܋x�b2��D��̽���4K��]��M`]�֛;~:Ǌ��:o2Ŀ4�f�H���NACo݋�t&���y��?v/#z�LU�[���c|�K�P�*#��C �6�ho�w��o>(��6PK�ۤn����t�)'w|LF*��P��*@�4T��+[�-���UTJ��N���qҝR��m���Y`��gxa�u&	!'�*��<�7(��6s�C�LL��E��L�א$Q�d�0�'7U�%8kI���P���7���]B&6Rf�.��̟-�~��]�#>������\կ�
��/ ]�c��|�Q}ҧ��D0=����T�-�n��)%��vz5�AY-���z�|mY>�b�m�NC>��q��X#��8�F�Sl�V��>�Q>�����)��ՠ���z�ٛ���,FI	>O񵓌��r_�+k�qK����XL_���ȑ���s	̄N+7)��]����쪳9 ��kp�A!&Z!uX����3^�v������e`C9Z���w��e�oa=��w��+�7�r!й�!	ǭ��&�k���1!FHM�9N"7v2���WO
w�S�N�K����g�B�t����	���?kHuK�!Ȃߝ_i�U�����k����gw �C���������O��9��X�np�?=��k��ۊ���	W��v�j{Zd�Qg�39:��Z��;|���x����Jj~��ѩ��U5�,��8���4nDk`�=�I��f��;�Wy�@5u�	~�y庐]89�MT����1k�|��TI`�� �K�K�̄ʪB
 �*���蚙�k�2Y�����3�#>p���.�Lۃ��MF����Ն�~��J�&NX\������H�2�f8�\e��F�;۔����}�op��I4U�%�/�܏���n��'�Cr��m�wK^c���`�.��5q�V*deTiϵFYKI��x�_q=���Bqc�͙Ȅ�Av���bg���vF-1�$�	ݬ���P����)MI	���``7�����\ݿ��J*^~�s�r��@B��r��G�����e���,*�%��	�륽�y�~����XL��evy%s�i وM��*o������D�"�͢K����3s����BK\��wyKm?�ʇ��ꪈ6ڈ�0�1i�/�*��n�t��Q>���x��ȿ�����ojۈ�T4 �)P�<Z�:M5{�?��Ҿ�H�z���m#��s�Xu375
�Ś��>��kl9b!��Mk��1!�3�$1�J�}�k5�(�$9	5�.��9�t����~�Kƀ�n�r�'�y?�����t��'ٯ���
���*]no��D%b��_Y��v�bM�o�'�[���G.�{,�BcB�e����ӂ�C�ݠN)>��-ԑv��h�O�j�h]�
�O��T)Qԓ��i���ܩ��k��IV�A�-��NZ��.�y��X�y�s�s ��3QI���s��
ZoOgk��X��Z��>2���l7Uph��M�݈��asF�3���8�¦A��q56(�T�ŉ�pr킲�(�'ٗu�!T�4�� �L�M+�4�*b��>g^b�<�8�
���ֻh�[[˽�R�<s��(J#MepfXm�\�;G��Q���x�L�+��ҥr��"�\ؙ7K¶k���HML�Z5��O!�C���5�8���2Y�����aw���>��[(�05�f�;�������n�;����I���a��z�s�4��7�`�h��B?�ɺ,+�2TyB@$v9�Fdj�X���Y�����e���L��q`@��Ϸ�̏ԟË���,�!A��zb.�~��d�L��������t��<�'#?�%�b��<���
t��B?�T��v�^� �����8��`�О����c:Z���!ng��Ju��ܭ6�� ����.�%���Y'�ĥ����)��"���d����?<�!������i��n�V��Q��Q�hD̽L8��[��W23�]��]�{}k�W
 ��|r(q2��6b�h�D=��9'^�L̸%uW�-�/�D���I�VA��E}ægR�$?.X�r���=���˧�F��D�$��ءJ��"����s6=�)����N���c�=o1Pq�����|A݉R��\b�� ����{�1{�{���7���m2e�h�-T�m����H��ZKLs�t�r7zh�I�÷��%�W�dp�BB������eÒD�}==��
K[n�ɽ�I�FzĬ�n\	���ɜ�m��Ǚ��,�4�T�7�Y�;^�K\�g�Ws�Q��F+�;��b�;���~�pغ�}_��c�x�����M���]eͼ�0{ب��GeD~㵂K�u���^�X5� 	A�G{�k�߶pSl#o��|m?u�*߻�F�`<JL��3�X�F�xń�#�"�#QJ���c� &�R��\�����-t�s�v��yy� h�)s��o��s�����K��]E'���QZ�����S���;f�����rO��N���'�.�K����F��Us�@��(42�P�[�|@i ��?r<��$�a6/W�Yq��.��n�O׃Jt]P�h�\���U�#���6
�Z ���{y!0�!�L$D���u�PL�;���&M�����ۇS��g�%�Z���������[ѧ>�0��t&�)v�z�sa.�1�⬚-.|c7o�t���S�#�O�m��]{~��6���u9!�7�6�̏L�E�Fi�o~Qx�q��q���8�%`>�o�w���u����8>�������W!�-��VH;�g�1�w,,�[p�����Ɋw�p���`����x��[���H�-�̡��ԓ$�V�b��䖍�O�R
QL��0`M������+3�ы���w��#�p�����Nq����<��&��Bp��O)�߾�Xy�O�u=s�����'V߂�{MmW��1��{3�d��	LXVC~�8Y}���o�F�>pwf|�hL��a�����L��]�X	��Y�Fy�{&K$c0��)�*s{~%���I���}�Aǎ=BnIc2���5��!\���{ږ%�=���-�5��ű�q���n��c�d�l��,����Lv����j��8�Y;[�/,��+�!���w��:ݚ'�8�X� ������d�ܼ���}�����>F%�M����{��L����5U�z�c�V>9�lV:�:�~��f���
�ZZ�&Lw)��1E`\�ml�~BeU -��Ϳ� �k�l|E�7��;���Z��t��~�x�0jj��#���d�-��̉��D=�=\���-к!�H�%���x.�D���`{���v�-���fְx�4�p��{խ��1�)���g�]����B����%��_"t�ǯ����\��[��?��O7����'?n������%9؁��E̗����Dv1A��!�Ӄ�چ��y�.w�h/}��U8�*�4͇T�ǌP��;�l]�t�Q�A�΁�H�$hoQ�0.z�gJ/��M`��S�w��Įxؐ��	�(B����Ȳ�\&�s���M�}[���93�i�L!���z�"�w23��wL���ٱ��e�s
&��+*{�������)(
T��+��'�>��8%w���O`�t��A)ף��K�s ��g�?����s�Z�������
?�4�E�A؍$&$��u��X"\�m�v���(���ã���1�D�9�{\�V��w�g�Aw�ㄜ��ܝ�ݿ洆]ϵK	K���B0Ws�W�N�4(gU�����[]^�j��h��l�W.'16}ǌ����ArLH�Md#�k	p���I��S�E�4��ͮ_Kn�cN;gN��?��\#(�Ƞ�����Ε�.����L��V��3����uYX�~CwBp���63.ˇ8[�g�q��=��I�eҶf�,\�	��n򶝩m�v~�)��ֵ0Y�ٙ�" ��&�H-�t���1���@�������Y�����M!
���#�`�L�)�ȥ��F��֦�8f@c2����RT4Z�sXp����؍�kRf�n�jH�7�l��p�ЋC�œG�-C^���Lq� MkwSީ��}\|��J��t��v��0�t�q�� :��w��������G�X�YW7#����?�wb]�a����j�����&O�b-Ͱ{��E�S���F�L��y�\-+�!�F/.��}�6�}OȾ�����Ji�٥�خ	�N�Q��~�~)�R���33�elI�w��UP���1�qw%���cF1�Y�7�`�Y��Ԋ�۞���� ��\�iu�TB�q��A�_��ў��}S�*7<��Jk� O���M���6JEam7ȼ�O��C�U����}��s{���'h����[���+���I3����w�N����!y>L�\1�4�~#C���� aW�,Y ��%B��� ����鉈y!��m2؝�7����t�����#�5M��]�2�Q>�?��EV4���ɓ�r0ɝ?���6 T<;�ߐa�5���Pi_�P�������֤�Q�o��nO!�c��ۣ��t���c��Lp�$��Y}��v�����Fu.o��F`V��[n1D��gU����^�h������i�߲s�/�~'A�����ᤲ�����	�(����F���n��朽�ßkk�w�Q�G,��������7���p�,�=��'��ݖ�ٸ��=N�bJ�����cHa><�HR
)��z=U^΅��j���z��� $B|a3FҵN`4�|��8O
]K�U���	�ܦ���Ų6�m�8U�&����Ŵ������|����:���[�������*�u�d>�$��.����=Ab�=,<�Q$�k�Vs��KY!��Z��`�=��=���>97���hB��u>�^c�����
�����A���0��$�8FxQ)�g�2�]��C�DV�y��c�(b>�[oU�|�7.�2�����@�G}�M����.aMYz�N
=�h�Tõ`�z�hz�\��\��~v�4L/ū�ΡrǑ0��'h�����
r��d5k��c��3�æ��7@�z�J�a@������i?���?Y��x���0�$�ފ��({"���e���f �ºNؙ_b���YT�C�!}������f�گ��S��w�#�2�3�2BUq������[��8�y���!�� 8���R�?�5�����Љy�o�!C�QM�0�k��o�+���3xI��,���qwM9����92�=I�$����L)����m�=����~��Zu��Afg	���N!�//�.��%&Σ���cd:^�dlfZH�����P�Ôv��s���pj���	�q��Y�q]��A�Eќ�/���f2�ʻ!��z!e�f"i]�[Ca�tC���ռ��И��x�)���!8&��}F�:~H�8�Ԯv9$?[�3#�andtz���OɎ{�����E����sB8
u�d�)uo��4� �>?�G�q�H򕢛��x�/��oe���(v�z�[��jz3c��,��.W&/�i�=v�Cҥ��%��g-ӫ��=C�C�{��raT����e �1��r���WF*��Y�Z�u��)���^M�+*8��$ۇ ��+��^��Mv��3O�������q0��{�6�;֍��y���bhgB���1>%|��l	�S|����Ϋ�u�uB�=e���sƺ�#���4Y�6�)��}�ϗeeu^�������$pk��/1�Rt���12�l�}������S �	�=�M	~鑭�����I�p]�u|YcUQփ-�$�� ��իK���WR\=hh�;FX[�����*ab����K9�ۮ[�U��	�Rh��]�:�F\�̐�S�Z������͵BpƉ����O5cr�c/;P�
�T��y��:uJ�_ʙ��!���#h�P���屣�}����!��/���{9y�2$��Z�|�;IѾ��ղ�m3}��ƶPB����~B�7�H�5+�{���%�N:�7��}����R�H�ϕ�ጴ	��pYo��>Y�i�Ҷ�p��,�А q�Sۣ�>����U��x��&�*�='�/詅r4�5-���JGY�I0@�{�+��Fi�`�!�&�5�D��'h^<uLz-|˸4��X�{��u&�x7�1�g@���/�Ț����BI��^���%-�g�t�۰¦����zW�"�e��Ո?,�a�9���{�gG1(�	�`J�%|S`���n&��e�i	ؤDaj����c� ��Ⱦ������g�*g�?;̈����CQs7���7�͓��N.�T���oK�*��(�-�>��i@��h��_����Ca�m�Ѩ�^��< ��ΐ	'Z���b���/�lN�v�KX7�I�ê��'M��4_�����c�-�&�jD���&�����#���r���h�J�v�mL"�)�7����k�.�'��9���O]�̳���Ne�T�v�X�S�@	��sx̸��)>�U�g�`w!���rҀ�|�n�v�u�����]��P��Wۤ楞~H�b{TMQ_���k�WN�.`��O��K�dqþ{p���
�혎�7�L���ã�^z��5���������Dn�Sk7��9��+���cʤ�]�	��-П�A3���):eɄ[/��C�}*��ԴETO��'I8B�4�PЛj)Ő���d�.K���̕N�s��֗�5�0�Ԅ>(�_����/ޅ�`Ĭ߻������[�P&��؈ 򽈘�.�7�sU���݅ ����ࠕ��2O5^���,0!��E�3)|g�o`IO
�O�S��6F=���9�/�o��csqU����Ǻ�h�" Ќ����n��:����3�̛Rp1� �QΔ�H�(?�;"�A6�z���g'7��30Y��l��Y�w�@q�x��if5C���@U�%��l���"Q�R�������i��W?r;�z���m
YjA��gr#�I"����k��+�Y<��gs��*i�Cc��F�ڎ%�ᶳ�~�8��,�X��\:��l���`&O���Ճ
Ö߅��BÁ	V�/|����15ԡ��i�����9ʡux����s~�}��0�b�U)y��6���SO�ڻ^�$OϮ�2��4!c��e�A��'*�F��D�E٢Al��F���\�'�D����Ub���C^>AXԅ��/��kJ?�m�`�@��.��z�F�6�[I�b�H?��$��MO>� ʢ���Q��m\l�9:(>�4d鴚'�m�K^���F1�q3*B��r�S��(����w�f{C�=���_�Z[Q�Q���"��Uq�$S�ό^i;-o�]����R-|#e�����Le�����(��.�����[(Y��䨵��n�x}�g:ŧO�>Kţ�����0uP*��=Ͼ��kF�Pe谀��W/M9'ſ�3Q\X�+�Cr;��*p�'t�Cq���_H�ؠ��R��Ճ�O53׋GG�0��7)�+�.\]��vWR~锳$��ݒ��Z��D�n���ϐ/�@�����_oA��$��1N�Q�peu��ˋ�����`�Xڂ�y"M�����-w���í|p����Cn��3s��\G!\L�ax�b���=I��BZ����_�X�L� �f<tK����;��oQ8T�FJ�$��Xn��VM�^/h�1:]P�dS�
���S��h V��O��f%�O�{�,�҅�	�*��;R�c4gV��Ȉb�42 �Z��4�+�|���;���R��B\Co�s!���OVKttoʸ�T^WN	��>Jm^1�6Ua��E��o9�N�%dj�~������0�TWB Hܾ��d)�>
D0c�V���ȖqG���,���.p��@X�x���E:�s++a��dh���ln-6�RA����: ~�㻠)��'��K��j�9�a
F�z3@� 2������Ö�<��x��V��!~�ǋ��ގ���%�!�P��3�8@���n[���c��Z� ���X�?U�o��� �������؍�d%��C,rë��w��X.�ǭƙ�z]��!# .����I=<��(Nl��9�.,aX$򚬫� �\�׍��\��򾯘�ӕ9�Ƅ�PϬ!lK4SPZ�e���z���XiDj��֝�n|Z"��.3�޿UK`R/VE;˒��ޝxrS ��ͫ��9.�lK]���_m���Zq��CL��GO�s���N^��wK(&ƈ��:D?t��6����e��*#�Y� �L���\�
Dg��6����Ĳb	 JR�X�����Sm"z��xHD�����J�ԇu�����܃*0�]�C&�'��3U��'��vLt�_���y-�@����)�D�/�{'�&1���݆_C����c�F{�1Bl�c����\:��;�@����V�*Tቶ'�V��{�U˷Jo�D�G?�^}c��~�(b!rh��ͅ�]Py��o���v�z�� ?������I����<�9t��7�����0В�V��I�X1���d��Π|b�����<��&��=���ǿ���T��w41:�6�v6(cER�RU�/<�����g�A�|1?������'_�竮pc�l���`�	���\>�cל r(�����(��M�0�:w�]!�C��$�Q�ы��5���قE�_@e��)]�z�68����Yڧg��2K_|!�:��}���+��'?��A��0�ߚ��*��U4<����8�TR;��B,3�7�'�-l���l&���#�/������h�B�i
�Wg��+-:�2�E��$�@u:��H!y���-�^*��xB�+�۠yP��
0��mR�'�Ӊ�VPSI��KK�X��@���z��UQ�}HV��W���n�Z�ٿG��|�c����Z;�hSy�]���s��ێ�]�QI`5�E�{��F���%+��� �2qOۤ�ɛMVv�w��h���V0��m���_��Jc��J�4=B�̙2a���6"	��_AsĹw����!~�E0�ث[�M"S
F
��_gK�G�[���gPCHÄ��
�(�8��c�m�����ϵ>�+����\FT�S���j_�h�2�{^�ؼ�B�j����6d����Ѳ>�n�t���SL�e��e��<� �i����U�{H��Ŵ����� 2d��N�b�w��Dy��(d��:�bF���|�[��w鿇(5�n4�D��X��ּ	TAʩ�v;7��!���pAGk���/j�;�x#���)����۹�[R�lc��S�^��A'�t��d��F�����4�e��%/�-HI�"��(��_�f�A��[:�7Wu���y�@��d�|}�(�A�W��jƫM���#@*�0��n6�x��@S��rApQ�zh @�s6�!�_���X�����?�e�0�Y�&�<�&��ԉRO%q���:��pKx���9ȯ͝|��̀nJȚ  ~ �,Q�����DܤK��qQ��;kJ�T�F8Y3]�6 �N�}qzi��n���G�,)ajL�2A+��N��������-�cՍ�6����%�{�*(�+��l�X�jF���<���L:���=�ECH�-��yx�jr�2��3�2t���G�3`�	 (t��7��\��X�n2���MB�tD�C��vB��[����I��I@޽���%g
�*ex6T��ޱ%;c�ق��?m��◶��oOHUm���7G0@�Z,.�/����h-�v�^�+x�k#��	�0`	2�Z ]l�g��N�0�2 �Nv��N已�E~��Ry�������
k$�!-�?7� �$��H$-iPJ�Bgx&ȴ�J1`�r�~�i���������h�N����8{��>;����
��/]qyئ;8ݏ�u5�v�x"�#�-]k}��J�� �A�.���A���=�ï�Xp'7���q,#�y� ǫ؅km�.�G߃�A-�w�K�_k'�	)��ͲƧrQFB��#P�?f4��V�9�xB���*�����S�ҁJ�2��6�mD |�y�Z�������ܑ�0Z)���,�#�.�+�+:�¡1v���y�s��-Y��[�͌c�$1���V��-/ �@���YM��{!�'x�z�*c�%
i\� 	����q�p3s�|����q��4R�hU�_�H��Q�i�q���\7*</�n��)���T[r��v�h�%�Y0���m[*�@��M��b��wg��fh���i�����Ǖ_j=�o2�\k�ӡ����K,�-����U��,���������V_�n�װѠ��Fq���P%7dDd��䘘e-����n�z��5"��Z��lʿp�2��Do�>j��1%ڰ)u$i�%�`�0#�]�
Z�w>��_��q��s��!�^�4���9~]�7�'�W������]���R�l�!~��HiK��#%.~�=o*��H��g��5oM��b[�:���k�Y���(��ffG�T�h1\�C�� �k��4Ծ
#��~� ��ܟ��-u �ۭR#�����Q�RJ�`FSk��d��&Z46�Ρ]��"��h6)��WH����K�w��X2A���aR���W�	G�-����� �2	�Ƙ���~�;��@���3�׾;|����߽tɡ���."10 O�����t���GԀq�81R�$D]�L?����KW�z#�R��4�[]���7/�"��c�s�{o�����5�a�=�*��|e�S���9wEN1�k���2���Ǒ2÷�oٹ��|BrL&?��տ:2?�����O�ַѽ�`(}�4gs�����AJ��T�_�����,-�y��x��ܚ#I�D���*Vv#O�X3��.2������ev�\�wMi�8r}\��3o�yo�!�R��%$�%�T��� �{�l#hH�en5+" xqg�=�ff	�A	՘_��y"���q�oIm�Lw���9� ��*��`����dY��Jm���R���M����4�A�DY*�ř��M� �<-���`ݪ2�%��'��t��%�j��x�{Pp1��<f�+�i8����F/)���Z��o���s�6fV�'<�p�|ļvO咒tK]�!A)~ϙ�]mIE���S��w)�L��P���sg�y� z�0���l�Ď�p6.r��B�s˃	!�+U
��\����|�cȠ~�O_��!;rw܋S�@���.����Y�}�<,�2R����	惥��Zu�-{lrd�y�m�	�m�.��J��oB
���V�Kq���{Da�|����F�#�s��3qI|-��Ӟ�١�Q��_����$��L���ok"C�x�h�ԛ�h�f	4aQ��sY6���3tP��0z^�k��%���~ejH���<�E<��L�_Y�IoY,�s���?,�(тs�-.̩�|�L���l�L1(N&fg��K^���Ja��9�b$����q.p�����+��z��] 16�X}t1'�M����Gqx���v�$f�ԉr��Y?�$��F(Nitٷ��^�"�{�g/������9Z����8h(.I5�R��	Vl=9@+t<F�)o�n�����ufI���*�o^YBhz��!Ṡ�r"啱����ʹ[8 ?Vz�Q�oDf��ή����{x�x�����J�]��s�H1�>;)�zkt�ٙr���ǖ�fOM:�F pp5�p�R�Y�h8\"ͅ�E�]�P��>g�s���; (5fA�{Q#���9��U��\NS�I%Ԁ���+~�����=j${�2ѹ��P`#�5��u.Z$�ve��޵V+��,�TTp�1b���<N�@��.��2%�x�no�ä���R��b�v�q�'��]�ae��O�YZ��Ǭ:�8+��,l0���\+-�_��*P�A���/��,U�:����=�C�Ca�\�&}RQ%q8���V�}$P�7�}hYTt�i�����4�)�SP�m:���k %y�Vx��̛��}���� �t���'W'��d2Ɖ�@�R�s�%AP�� \�l���V$��ʚ2>_�f�k>	�,�.y���y:�6"�^�xD���Z�B�p�ᥥ���o=z�Ǜa��	|@��D�|���n�y.v������^1J�_0�1_��r���"$����w��6�at-0D�C�/�ڇ&�K)���� Ѩ�n���u>��N`��0��(�'�I�!Y�fz(�-�S���몏�r�O��䝉
����Z�`�}X������e��q��h�谹�!�fMP���{�:���A)PsT+����C$ v�]�k�0���M5{�E�u��##V��H�	���T�B�g ?w��0x3��KwB���-���0���ȴ�#�� ��ن��F\	����:����� ��O���H-z����w��]�	�k�}��a����6�":u�z!/Q��(=�DI�|!����θ��7�e�X��14����,�p��`�U�&�^$I<4�*��
�m�6�G����5pV"k�T:l�/D.����2F�XTU�;��E�\�d�'�?Y�Ey��V�{郑\T_ꚔyQ/�G�(�$-��	��&!s��|���`��c�vo��0~��n�7Kdg����6�(�?�� ,2�$����4���{�&�@�z���H�]"a���q���k ���*L����"S��P|�d��V�mg�\�\�X(��#Vz����ܶ�]��)��;��=�e犯+��A@B8d�2]I�-p]̔� @�<�y�\hV�@>��E�x*[�� .kFYS�.�Q|����v��P��fy�j���H=
Q���\*Np,���n�s�3��MԂ���O�(�|����@�cG���Y�M����Y�:
u��E�{1!Ԝ]���*� ��>�V̱y��y��*f�|��.�Q�и�hv���Ƀ�w9=���s��{@�f<v����6��M�2{��t��J9��ZỼg�<Z�]>z'w���C���	x��|F1� ��{�g�a�b�agaDc袎�̚j��0��O��h�֡η�PJd k��ds��VS֢wY�p�.�*V5�`1����*���q-8U �h�4y�ϖ��Ȳ���t��4'�j��f*��PMm�dqC;���\���[���Gl�G��:����٦d|�3pS4��XM#��ŕ�`z�2��)� �dōuㆪ6z*sf+�mh�$�%|q���%�~UB��vn`����,�Ѡ!,�nK�����5�]-f�{�v/�o���$~����,�$�Y/�����>��#n+ʹ��X\^���\Vw�T��~�t0�M%�U3��['<-���;/�W��5g
����LVa%�G���K�CJC����#��l�� 'Wc���au-ς��2�Y4l�x�p�$���MK%�G�F���8�tXgY�Bf�g�	@�b�8R��lt�êF����ОS�$�,����~4�L���f܀`,N���QM�zM�����S�xAҿ���\�:H�CgH�$���Rfl�h�-�\U���.f�[�8�,�=o�vvt�}X�6J�ݛ�?��IeWh�HP�U��}Na��DZ�w���u�W
>"|ϧ�b�yԼ�&�$c��K���́��S/X'k�I��ѽ02�sT��)4�
�������΂�@F�(G�n�[���*�/kE�����w�ۂ6�4��+���3e�IS�X�4�0?K�eX�voS~�����{��+��r�nDF#���@����ܛd��%C�� �֪awW�����=�95I�B��{��?�R��~�+H�k_�f����^����KF�^#>��V�\Z��Y*\2�O�L��{�<p�0>>���h���x�os�����|�k��܋}fmmS�
��X$�)��#$j�|zR/`8�r�$�O$���d2���x?���-��@y���-��|�l_j6ж"^M��xQ^��@�Y�_F5�G�s��;�惗��L��������e-�Db�(59�e���KA�	��U`	4`A����,�U �K����{U&��9$킗�e�dI�}>���L�{na���	n�:�VtW�N��ym��𻂧/���G+q���rP""�f-Gj,��6���sp0j�b���&>�m��%a�n�.��2A4�%#d�s�:~8 ��ۃwy��*��x���(���krw�1.nRG�@����~ �D��9���t�7*���L���P�"�g�<�l%��ك�-�eIhfZ��Iڧ�׭�h����/d|���C��hk*�p�T$�հ@�C���]j����պǛZ��F�r�}��}z�)ڐo�8�7��(r���U!�dߘ_N����g'M`_?@�bh%��	x��i0�fu���5��W�x>�|��ѓ��Q�&-+xp!���e���>WRh2��o(p�WUG.<��'� ���)k�ҁt1a��7
�G���]F�ٕ����]ia��@�q�cE��D�F���W����\�p����D-�fBc�a`c<�� �t��_}���eE'��j��T��d1E��*Q����Ό��5z�X��=���c4�m`�.������Oߕ� �^
�*E�ߑ�@5�L����5��v[�^���L$I�T��Ǩ.I��RaY�67#'�9|D
X;+�ⰃC� Ԍ�g�He�m���?-`���Ibr��s���t�?�����;;�W��&�'I#=v̪k��N�sȷ�}~�v:P*?�Q��r����N�u�Eϣ��|��	�q�}/*B9r��}a45��.8�GoT�0�"m���H��c��{4T_�l������9�O�ujh%T�	�F��%gL���4���l"�� ��i&s���$�ɳ6l���Pښ��bw�	�'׺��g��_�����K�qJ}K�
��+wg�1#�|I����a����i�߰�jD�q����'
4�c#�Tk�w�~�r"G���#�(/f��SU�O��A����B�a�D��7(> Fѥx_n����^�(�*��5������ֱ���z+��-w|3��E�@��k$G������c�_+p05No)<^9m�66pZ�bX��>2�j��'���i�8z�oZ[
�n��_���YYх��(惹.D��Y:5$��XTq(�ɽ�s0�"x�_��,N�(WԂ>��\_�����;�Ӑ2�&S�'ѻ{_Ʌ���^R=M�k��N��}ٲ�IT��s_���&|!���zt��ʕg��c�����g񄤦ãk��	��>������pRQ�`!NQP��H��r�EG��ՠwT�_Eb&Gh�T"�`�&m����C�%Ue��x�̳���j�g`H'")Ph���jӞ�:b�pg�h��ݖ�9��P䱧�[_2\Lθ�xg1���b0��N �S��l�@Y�q�����X ����IDWr�*�����?)O�z���Z"˅ۓ�g��}��%�u!�U
�_�N �M�P�7�[vzr����CO�+l�(�IbK5-��<]\��c�w�?>Z��>	YF�çD��Ҽ�7!7X	�(�M��w	�*���~��J)w��:�٭Ae�Z/�� ��+�%���mF���h@�㔬ދ�?i�q�N8d��(�:��ժ�h��!t󶣔�����Q��� P���6y�#��M���ؖÏ��ᯀ�~��[�(��j�V�ZJ�y��*��j@;��>�o4��Au�۟&��Ri�G���&��z�4���q3��9^^�ւ�ȯ0��&cϮR�]�ήb(po��jE�1�g�e�����uu����ә��lV]^���1���!�������*���%]��v_7��v�6o�T�>�ʟ�)��=�m8'B_ܽ��K�uoW~bǛE/r'̔�V/ j�x�=��@ϔo���r)���e�ZY $K�3'�	`�v���橪���GC���,V���|R�/x_r�n�@q�;��T��x@",Fl���Ua9S���������ѓ�y�m��a��/,R�qҖ�K������j��[!����<U'�E��[���^��e%�ܛ�[�O�> |��0)H!��p��G��!z�{�z=}�߭V�����j��	�s�]���"�21<�5�����K�O�zg�K����S{˴OZ�u���=�?��`�b�YlO�8�������8^J	��2:���o:]��WHF6���ً�ep4�rcY��I��>�i�x���4�g��v��H4��Z�-
�W��BL<v#5�x�JG��w��~o��w'�i�2�>l��/���g�x6@�PL�d�����T�e�Q7D�Q�Jk��)E�h�g�a��O�s�������>�LJN��k�H���a�3wՆ��ۯ[sV�\�Yz�t����AG�̄_#bk����c9C���V�Ii�T;��?.�L_3.�4���?�]R��߭��ϧ>d���?�]��6��RMUT\����I湚FYb�L��r�h�ٳ48&���)�=�,Z�-�����*�h6�
�ܛ�Q{�dk�����֧����
^пt�@�e[�4E��.Fi�1� �9*vk[���g��MG�S7�����Fg�\���4����/i�&��@&��YV��6X�/�߀K.����ͫZ'���xq����	��6r=A;�Q����=l��U	g��wP�9S��yi�t�p�����'��
��r��k%dDo
��1&��o90�`[Aʃ3l��5�W%�����)���
���I}#�j��(�-6	�m�2D4�z`���guQ�ElM��'Wj�ׅ)�K������&Fə�(���Pyy�������o��.��C�����K�ȉ��9z�&[��YT��ͨ�P��Tvݜ�k�Ä)��3I�MŮ=<����5�K�Bt��BRj+TedՖչVxq�8͆�`�5U���w��=Z=W����ɪS*�lAu�%U�E��s�!f#�G�*�v� �ڡ����L��i�w3�tRح�X�o� �a��?,���',8�
,Q��'H�ݺ)���Q�	�I�	Y�Sm���<����b� -��b�'~5���&	O��gI�#��*f.qSl�>�X!F��(�N�5lQ�cHM�3KD���)����"�{+�_�"pGԼ��ͷ�%�m����iFy������R&5�G����=��h���~N���d7؋��
2���%�H���4
iY<��]0�|u��MZN���C4��2t3���@PX�i�ɱ[�g�W�-A�3���3�O�ݣ�ڥA?e|�2v�V��� "AC�iʛ�sG�D��EܹE���'{8l��1���S���{t��)+I$&l.�Al��F����mRˡ˦"� 60ʢg[�+���5@�` ��`�B'���C	�]@���4 /�>����w���pR垌X��BzfjOA�T���=�2^&eԎEۿ Ĵ�2Άb�v�~<S�XMP^4 )���#��g�z!a�k3����_�w��nC�)�qCВ�ذ�/��-�i�7c���
����I�`�V(��~Aݳ�[R�D��1۳E온c��/`�#�2�0��I�PC����nL������):>��(�Q��"5&���eª�빡@$�Q�4��W�YLCV	̐��٪|��zӒZ>��ʟ�D��|�?��u��<���f�|�B����k���Y�j�(Q��ū�n���أ���L��(������ᚮ�LVb�l5�u��ۺB]|��/&�>Z0���v�׀�0���+mל:4��c�8֭�҈�٩��)y�c\��X2�9�{fyŌ��:�K�m{�pv��iYcb�C�4�F_+�����T=�N�'�2n�b)��k��E�zL�8)ܞp��.�ZM��*�WWT����C�~Xq�t��z��ns�����o��Mc��"s�d{�pE�8�}�����ݮ�M���w�,�n�%�օ��X&LE�|���n��L~m��G0���fݔ���9����I�7���4�p�+>�!@I��PT��Mm�q��Uq���R�^��5�ۿb6�枹"'9k�v�s���Ek�ǤD�!�|�o��G�P�g[>��E2��}��v᳊�P�c�QA�zh��M��\�$�pc�6a�
ط�wJS��I`:�$�ݫ2�/�l����,W���p<e9�>4�)`_^t�yh�kn,��r�`X~��U%�)��G���-��H��N}薢nyx+�Ou��N�?�e�E�d�&2�A/�v�cM"�>��Bopa�R.!�5w�g�zi�oD��-diݦ��(w8��>����P�c}H0�'.�ߟ������&��H���6�"�N��b@�7nAd�Z�@>V����8�9�X��ZV0ߗ�QeR�*FK�Px�E�}"�>�%1��-�i���W�n+"9��F�8C�~���{8ޜWlMd�:F���c���V�Z$N/V�	3	���'�6X�JB0c��Ձ[�`��ܜ��:LK���J��ї���G� O���j�Y�ݴ��#i�q����-*i�u����(�ջ�RN�)��m"�xN��Bt���P����d7�����S�t��hژ��Y�[�}�E���G3l�/l\�nUƽ!Zz�� �tF~��t~�����Q,:��m��j�#���,�^�foYZ����7��a�#}]�U
�n�PY�jZ�<�D�T<�cή�;c˼-��U��2�8P�����B�����sO���2n���	H�!��Z~��t���o�?"�y}_r��0S_�#_�+��OY��|�+�<s�|�]I�h�ԝ�"UT�}��@GS�D}kk�}�^1BG �=��-S�2��V���m<�g��f�Y��طGH�"5_#�I�<PC�P�m�&n�ߚ�T�/��gu��h�2\@w�r�X�d�bR���p$N��ˑ�����Q�<������3���VW<H@³~^h>����("�zm?.h�8^  ���l�&�͉`��`[��C�L�DB#t����5��0�H�?��"�`̯kR.�݃9t�`Z�r�'$����}�)�>p����B\Hr�0p���pY �5�z�T�7,�v����&x�iם��h_�-l��) �����|TJmҲ�Ȼ�ܲ?!}*
��9ʵGR��2J���V:/�}(��ъD��{�X/��V�.�l'(q���(�~��l��WƢ��D�$}�M�� y5~��9u����w�G<�g㓲F��L�oI�y P�]�Ғ�Ba�$���vm�*{>��c}c�W
�+�-x�SW�y��c��T��C�v�&S�<�8�qC�o~B������@n��9h&��b���s[яB��@�T�IӔ$�Mʩ��m�V�H ��6c������۪�!.l|�Tt��Nx��`��PbN=��r�ߏ.L(���BԀ�GYi���?���0�龁gRL�k���)���S�G�[P�$"*@EP�XG��5R���nB� /D)��E��Ȕ�c�V�m.v��[L�9P.َvdT\�g?��{4�Tr�EW�r����~q-;��q6<������>�w�e} �q3&BM��8�ꆂ�`Ry����ߍ�mxO��� Y��0��ͱ�.^�	�IAN��!���W��+ ��Z����h���A���Z[��6��ո�o�-]lpԉ�����?Cwl<Nwh�2�+	��1�9` �6�o�r+Tk'*v���%�P�
�xEix�HۺV�$�)���<�t%�� �c�
�EH-(
��n�0�]�!�#�a��2��#���� {n��/l;�^ؚjpل�	pU6ب�� !�n	�zL0��p9�z2��=w:�X��/(M��6��g�/�t����U�E9lr��B�^l�[<�E2h�Ζ�֡Lǅ�T	iޯ�����'��xz�-NO�-p^�\��XJڞ�|V�8��4��6Ə��Ӱ��%@76��Cd1�eF���~�Q��<1.:< ��'XS[�M��D!	pY��7&�� VK}�v��V$���)�6��{��_Ռ�i�Қ�	�p�CF?حR}����bTI^�X?����A[;��ą8!�6�Ų
��3�S�.��f�+f��d�
ˋJ������[e���UX�- ����ws���o2�yҞ�*hbt��Ū�?��=�d7H��|�"�[Q�0�W7G � |�#�o�>b#�"U#��Jk�4��iY�d޾Edm��-!�`�Q[O�� ф,� ԰E��h�į	��V�D�)�)̯�������B�;i�uX�s!T���,�~�����ߵ[ҋ5����vϞ>��@(�O�����hqC`���o7�Sw�Ӝi3�䝱�,KR�ڌ�?���F1�d|��������G�N��%�,��<D��P4aF��^�\����XM�+�ܷ���o����E5�8?׌�G2��6eƤ;�ߨth�|�3��x��� �q�I���2mEh�A��t�a\_I�
7o�=K#��#c��@��qk�K�/�(�5H�ĵs�*%���C~�M@�7�\��Q���aD��}��S�VH�'�x���Z`���:�yB1]�S�O��F?��N˪�3seߢ[��)ñ��3��m�S59��p83�f}~j&�h=:8([�_�@��n���g����O�����0�[�d|m�S#.	����m��D�8L��b���_j	���*����?��"3�r&��O�Wg*��l}ȥ��fD^K6��mm N���Ga��6�V^�bMLjYd�w����#�x�gbvvSgS�Az��Q�gP�c�d+
�XH
���_�c���Pn��!��߿e�����Rw��8��5d!U�O#�Oa$�o"wY�战�(�#�ufn�]�j���c�^�WLVK������ݔ�<��4?Td{�u�N,H�8>NЌx���|c���,��Ћ-?Xh)���do����L�
՗��'�`;���jCIUvD���q�e9Z�P���hn���Eu����:�k�����!�{�U�u�.��3��>�cK�ܹ2�ͯ��p6+l�x��$\ƍu} �c��:0�ͤD��Tj
�)t�+,����v]~Y�>n�]���g���!���L�z��=�ZHk��d~�2wJ�1���a���ڡ̗�%y+2)� T�Xid�]W>O� �������|�q��������
�Q��g�)�*���<�d+���80W�uѳ����"�ȳ��o2@"HB��{�L��GE\����W,U��L��Ԙ$���if��p�+��F���`�s����q�וS#u�yϋ���K��Em���#�P���q �1#�rm�	w�Nu�zzS��Y�&`+y`�n���L���������{�պ r��[�̢�q���i��P$s�h4T��kOa����|Ђ��=_&f4��n���a�����K/o�c�W��+"c=�� �����SR��
��m�����8 ��I�y��������R��cF��$Y���<�. #7 ^ 52�r2Ӝ� ��^'ʛ
\�?�U�x\h�7�ÔS����U��G��'�}�-������QK��K�<>$Q0!>J�2̨���`���Z�9ڎ�,:T)�㘶�L,ED�7Đ�	�,TXn5O'����T>�k��:֕ֈ)�<8�u!]��5��F�(F�u�(a��J�GW���/A�,�AQ]��M�;�.O�7A�ӳɋ5)��eO�/Q��?�d7��u1P� u�
i[4���LK�n��ȧ��sfe�N�ɗ0��9�����?�"����S���I,�%�-�0
��g2X���j�l��b��{71�x����>�����xF��oϬ���3C�\V!
v�8"G���HŭIo_�m6�ahQ���@`���II�GlQ�6 ��][��	������S��������0����Pg'�M�]*=e��bmPN��>X[���#I����]���$Q��O@��k3��p�
�Ӄ�L��k�G�N�펯����Q�m����,���d+��s#�����=�M���XV|���ֹ7A�l�������V-6�rh���+��E�z΄z�&6��\2�Dc�_0\���l9���ys����^�T�?pjU�ɿA�-�����;�,�����Ҭg}�:�[��'��/�͉Kh�o�&]���wm)�?숸�O���������-t�M @�|�+5��v/H}��{ބ �|߻H4��r�� �pq�Ҵ�*��H��JO\�R_\]F������	��S�.�^�Å�������� fɦ���7KwO�Qdz��u�$?��M ��rQi��8�l��:Ŗ9�_T�|�{�̦\'�袅���gb��G7o�'�ph�QЏ�eY�z��y	���;L<$�/�*X����jt%�Зz�W�| ������5�o�.�̻{�g�ތ�F��()	�,B���J�8�Cۼ���.0��i>T��Ԇ�k�$4锱d��3d�h�RA��T5l�,��`������h�}]5Mw���$��uZ*�?��#���f����Gl���7��m@�h��x�N/{d��'��=��<?/�R41�h�P�zòA�b
��X2Tn���0�xB��>���E ���>�l�oO�)�Y	�<yo!7I����W�Gr'd|-�	V�s�g/A�T�j�D#��<w����HM�K;Z����@��I�mmO+d[��:�~��@����1�e�7���J=b8�o4&��õ�	����݂�L��;�u	�˔�ur{���"�k��?J �u�J�0?|=ro|��׏����9�wgA�#���ک��V߱��~e~P�
�O�B}^���h����i�T ��H��]t���G���I��R�ks)���4���z�2�k[�$3��^���%΢K������U��S� ��	�7�D����1����F��)�$t��>��V=�l\�hk~V�kX�|�0��t!�9�n_XƜ�B&�/!<H-B�y
-��
��:��QB��k~y������Uy��6�^ͺI��u�$���� /r�z�Ύ����/`�ࢇ��uw!��Xy��t��eH�N|�Lܼ�yA�K�&U �Y
3�[���'���Y�&<�l:i�8z�<�l���:4��>0N+�!\vT�FxK�u�|�$�e��3��������?��&���#l/��G�:btk����H���Mt#�ۉE�/�G��N��LP�5����%�xɞ����Z��t����F�\z�g�5�� p���o��h�>YO���Ó]��E�R�����G�H��<9�qk�����AO�c>÷3�ח���`3DڊM���.`�G@{�.^�i���;�e4"0%h�)9�S
m�K,4����$�`D�`��ұ#%�Q������l;-�{0x���6���?�MCH�jFh��\Z�n /�Q?V+��<�z�d:��������)�Ǣ�0
��[��;�bܳl<�jYɿ�C�b�a"��R?~E� �d�V�P4WĞ`��lE^����C=�eP ��ν�5�E T��� 8�P����]��rADR�"d����Q|��|��+m���ť� !YP��D2�DA�ċ�_�q�,�3�G�1JE|���q[���I�=�3������Ђ��X�#���:�۪�l �����"譔Q,�~�v��fCa�	'ϱ�?�"���"U�����
��k,�$1(ԙx&��\�Z��u]�%qE��șm�(���Kz/�	K��k���!���[(�*�#Ukpc�I�r(��L�zZpR�Q�A
t��L��/������`�b�e.Ȍ	PIo�3�?�:_ s8Ǡ�S`��/;����W��Zpy�F���D�V*��P��/-�ŵ����:2pgR�q�b���j�0X��ΘM�0P� �%^�0h!瞍 V��r�ꛦێ�������n[��VZ��@��O ����I"�f�h
2��w���u*9���b:�8���V0P�F��K�*���X���W�]��A���	�PS`[�R�x��:T9?x�x����8V�;��w0�nH�q�ˍW#h�#J��r�0��p�3�?��V^�,ɛ��{E���I0��r�P7�m��Ui{d`CY�����O��1M.��"�qe+���I.���AwF�գ0
��7!��)ր�-��Ѕ#G>v2m��[2�7�p����67�7j}�(�����S�tV��1�M�e6����ٰW*%��n��Ѳe3,U�AǬ�l��V��^	.�<�`�V��n��b���2�i�eG�������Sӥ{$l&i�G�@�c���w �m,;��J�|�q~�9�7)j�p��{ƅ���	?Q���r�
�ē����'�B-���>4G\�ٵ�U�K�?�����!�Up8��3|��[P��:�c��ԵM9��b��8�xŶ��_�l�Mof4�����.���;�R�K�Y?Rk1Xf�oPÂq���Ie�c��2�sG���-��r.	���E][��S�{�:�Ve�����Ҫ�tj��=N�������5�G\]��.�4Ͻ�Ё�@GP���䱣=�"�"���3��}TQ&S�z�Vq���D�8u�"˱�w!���6��g.x�:U�3�ո�i����_��2��X��E�|&�3��Ck[� ,�S�ɹ�[;T貨�1u�0eU#�6q]TH���(I�z.�/q�;cɧ�"�tV�S�pA!�{D�*	/����]@f
�r���J+��'�t��.��n�?���PSP,�ɺqWk`?x����&��Z3Bo/�jI�K�J��^qu�i� %��bD2��B�[��oi�!֟#^��"��(m!�@���/��J��<�����9�}U���MN��U�ɭ�d�"b��e
���d�F�Eu�3�2J�2�|�cG��΄���VY����Hj��M�Qe3B趐���}&3MJ?`�L4J��ƱT*v�;)���l�ёɽWު�0[/��G���<�v#r��>7! �d輦�9z.�%���!��[�~�����֖��҉bh�D��D�;T<� �"ҫ���1!�ח���p�Ad� ,7g���J����qPv#[��j=+5D��3};T�+�/dLi)�`@��T�z%/\g俜-nVstJIR�(���nt/�eһ�XԭF����6�.�\t��� 8t�?�g�%����c�`�h
�y�9���5kOw�Qs���*0���:����Qlx�����n\���7�DSҥ��>�H�O�Y^1�%ۃW�|���j�nRś\VjM�=8h����oyD�V&PJZ�4I��:�.f��_�6��X��)��.X��We��}{�Abi��X���{Λ2����x�'x��ʫ�)��K���;_�3	���5�a9'�1�����Wݿ�)sǐ���T��X-b�o�(P�sу���s	g�P%/�7�����|�[E�(�G[(�"f�"!-�"Dz��?��H>��L���-G����B�T��|�������7r�Zbz���K��Sj%#fM%>V�.��5-´��-+ݵN���O���+t�
�:B������#�;}�m��M��ȳ���E5aWh�\_@ ��t��ɓ>�g��#��:��b�!�'��PR�sTX�x8~�6�o9Ǳ�I�k��s��v
�t1.�8R�(]0Æ�OE?@�#�AL!C�\��=�aH?�s�k�%)��}!o�*�@:���V�Ri�uH1<��~�C��� %�]�����i�-.�C�b��B��[���PH��tF`@��!	'lu����2�978TL��_!��A��j3m<�j�)Z��c0K?�{f��<�3�k��u�`� ��D?���R��q5�~���(2-M ��{q1��1���=�L�i������
����K�I%�y��7����a���]��̸��0 �F���,�s/`������h�{��@��܉,~��U�&~�$0twZ�R��!��y��
E
:�B������c�4�T��9�l�mO���*s'f��"+J(D¼?K���D� �E<O����b��lC�킽�4�	�ߛ�Í�����;��jo+Y�޻�i�>]?����}V���S����t���.�|es�bQaP�,ı�?�����5}�f0���$F-q[�T��dޒ��<j��$������������1y���uD��I�{���z�2�`� xϢ�g��o1�@��4ԪJh`.fB��'(���.̍��0>0��U�6��lkk�pY��[v��yS�qj*�xBz�hN�*p�&Ҁ�A���uHʏA�]h�_4@U�d��nٺ�7�g��\��\�ϱIA_�4�	��k�?G��Y��L:H���.�}L�D*��`ª�F����7�N�>$'M�h0�i3	8�5�>)��d)�7�=�t���B.�Ū�a��C)���2$k��iR/�Z���Z��������s#�A�w*��zav�_���g�����v���;x�_o�q�ے>i:N%��F567���Y]c�
9ڑ��ZFqG���;���U+m�̃��o�B��($�YᆤKS�:����MU��J��4>cBT�jp��#�i ��t|�x�cH:^B/��<.��j��'Tw7-{&�p�W<�#���ێ��݊S�+�Ծ �]�S�$�Ԗy�D���}Av���h�y�z�S�i�Id���!��N�n�}�HL/�}�j����Wa�g��+�y?ݓ��-Z���w�1}�.7|��z��t�ŷ�B������� ��<f䐕E�� �W���S�b�e�����t��p��,�S��*�L�01o?��XFIK��Mf���$LS�C"/��&S1��q,�,�ڥ���Z'<e�GqX���L�%�'�<��jH�����'D��5�J0��H˪U�zw��s,D���x��,J멍��U�Y���tË���M]R��i�������Kx�3�JJaC*��#�a���L�O��o5���%�lq��}�V�X��E�q�G�<�҆F���Xĉt=(��5�틈	�J����A*�*JB��	3�N���Bb���kԮ�,;%Q\��������4T>4��˾8{%^�/��q;�Uu�w�9~���[�1�v�K�Uq�B�Zx�ٮD�##��p4�T��z�eI��?ݴ�j�IZ�W+��^y? �F��0�Öo[�jCLWcg����p�!�Mi�x4s��k�$7[p��܆�=侦:�/#t��b����#;�D�Zr.(������l�pPԭ�]j��D䙍�c dgg̡V�{m�������=�^ɾel�����> ���'+����(��Z?�X�Yk�l%�����Jq�
D�²f����S���Z�'��s�;����0�}�"k�0ܝ�S[$7�z`+�ݢ�T�,�+�N6�`��+#�*�|�;Y|���
��|JR�hq�[���Ap��ϑ�<)�"�:�y��iqɚJ(eQ�Q�K�ǰv�h3���'G
��g�	VƵ+�fv�Z��,��Y���V:j��hdU�S��+�S�ɌH�eRv���O��8!lJ�H�EW���v��a�reyP�I��Nu���ã�iْV3�;P��5�1���'�C���j���p?)ɟ����|R�|��,�rj��:���o%>	$�2 hgˣ��c��6A6���[+��h��့�n�'D�8i��^+�
�+���l��I[����[�?���3 U�QLF�u�h��wn�W9���f����|��_ּ���&]�(?ǵ�ޞd���V���ᄢJ�,UuA҅Gm�������bZ��%JWU�>�6;1�5�mv^Pr࠳G�m�V�U�����+$E�3�d0F�R�g�!��!0��V`�zxv����_r=�n�q��'b��C��!#���_����x�Q�k�6�q�:0�x�[�K�8m(V�T�������m�H�Z�`�oy\���G�S�<� Q�M���H�Oy'���n�+�i�g� ������vX]S��q��(B_���Q��zmŇ�]�&�X�D���J-�O���5�#㥲�ތ�S16�Uf�'��D�և֣f_U�p�Q���q���; �/��ў�)�ͧ}<߯�|��b��o��v
��Q6� G�����dYZc�Ob�N��0�����^`�)���H0*��C��s�Pp�9sL�0L��Ċk���T	���%��5X. (㒌̜@��"���d�X�<nݦ>��[[�R�f!�T�F�����1�g�1��Ev1�!��-��מ8�l��1:G�^X(q�9t���SElPٮ����j�N�b<��D͆��&D�j��wU�K��N�SB錃h��Z����P<��b,�2d�҂�!��'���(.��(;�.�Y/gR���|�ﱸ��kUi��:�x PR��=K���ZY���s6N榤�f�H��\��&(��N��+F����-��B���D?m�\y�H2_L��>BظXd��6��6�b4x�w
����V�9B����������ș~�u)n;�xf1�:t?X�e��	>���f�d4]��a?=�P�$��q���?]e�j�~	�=��L�M��}���ܨȓ�+eI�sņry2?|�t���U"�xk���7�����$pz4�\h'<J��r�9ТS��瑾.rbc�܉JE,
�pJ�Y�_8( ����p��؂A
�=�wJw�Ѕ\���?��╵��i^��ԋ��=��RQ��%+;wQ�����L*D�`��Y����@Ω��l�	���1���^�&uQ�X�tA���HO*�
Y纗�zE{/��~��֣Zp�8`�L�A�"�4HTLA��ۥآɨ��g��[�u�����X̗,n���Z�����+id�O�W���\?%��a�9�-��s���W�@���n�q��0.x�I[��[���0�����p�6}�ȔXV�6%x���-?�k�F�����ߗ�t���ML|[}��*��^p��F�ِPh��s}�㘴�OJ�%��B�9��m9���1%hĹx8�7R�R�d���;3a_Ě��+[)�G�&�fNc�{��H�rY��������o �y���[ɝ9w�OgU�'�_c ����śr�mΒ��{�� �։f�f�a~�s)X�S�,�P�`yo��S:���z
m�Bv��d)}�X��L�:�����O}r��O�\�X�=n�m��k��3jyc�^,s�x�����AG
���35s�m�O{���������-�@?���A`,���D�<<�i������սb�A��ג:G�Y8sW��뱅�:'!��C���mF��O��\!�mS���fU���71��OnXm�����gkv^�׭W�&���p$��}~s�l) ���\	+T�c��FA%���z�I��P�u�I���[�79tϾJgɊ`, �aX��*�Jt6U޴c�xBz��aVQea�����.����j���&�I;�6gh���H�C�l�M��t,���4�+���Cv[����P �#P�u��R��ݐ�0}�8z�^��@�!�(��`ޡ��M��Qy�H�A9�A�KG�u�N�L�0V������H/
"�!P�Ac��b��(�|�^8�<%DI���$P��o��	��[g]�����4������Q~�����!\�iT����S�}u^-~`ʙt��
���A^4���"0�=��(wec�PRm�h��C���ѣ�g�L�w9�c퉘I9���2d�'�F3k�FPc�����w���"?�;=���}S�=<A�~,\�/\	Q�6�cvF��Rv�;P�=�e,ь��%�����%E`��e�ɽU��o5ݤ��W$'.Z��^��.�wbPP�W����1;kj���R���b8})����{C{�����a��[O �B�<>��~�u.J ��J��н�q�	��16:�Z�ǿ�s��6�]lԓ>�M[����-�6x�*����i�6���?��qGvjzz���"W'y�'%ݱ�_�TK>t6�:_��g,����2;��fq���%�%�G�2�a���T5+~!��=�r�����6�}ʌ�!չ������
}}�y�j� �
�\�_���rcI���N���A���^���������f�P�ܒ��DIR7�Sx 3:�C��w�����k'g�>Z�XE����j�
�wMG�O��NT*=�C;�N_M��L'_�J�M�2�+`�#�q�ۗ�N�[��m�ɭ�C�|~���=yj���f'<���ŰW4�(��2=���,e�gk�XsӋ�G���Y_v���	#������n^2���d3'2���i�kVl�(�R{��ȔFq���	��� ���}����%T&���y�99��!I�h�q��0�ƭ��IQhvL*�~M��+�פw��;ʺ]/�w~�Ècp_~$��y<E#\s�#�׌e9��\��V�/�%����B��y?E�ٛ�HJxAY���8d�����Ŕ��f!4��������H�h<�[��ފ��8�E]9�+��'J;�{�`�Nd-�s�s�2>�;
������S3�-4�`x2�3^v���w-u����S)mj��h�Z2�T��������nn�q7mf����*�X}υl{�����BT!q{z�I6����ݮ��Q9%md`DO�ᇍ(*I�Ч*)8j+q���L�����df9~9����7,�9Pt�;5��k�Z2C�K�!�O�|�R�Y���@�U���I�@�l_�A�ma|馕g��9��.����4�@�ĸO;	��'����1^�����u�_z�:�	I��3�ݣd�p�#)��Ƴ�:`��~�wB���}��?�kO�R���N��\_He�^��>�fdQըWc��羯^>0A	y�y|�N�0)���0�Y���L^Y��k�68��%qDE~�akB�4VHQO@�F?�1Z�6�됤���lt�".��;�-b�b����t��p_�8��u��RY����td<�=��4��~�|[��.�˫"2�B����oXř}�K0�/����N}@1.1.��l�H��#�.!�W���F�	N�h�tj��c!:�Pm��8�h��W���YEъP1
/'E��5b�����P��D�і�Ｑ@�]Z��m�X�Bܟ F�`��=f��,���lM�n10Krsؗp�š�t�U���p�m�n��<����Ge�Y�.�ЏC�
��ʸ�.��<�P��,�����Dd� !�f�\v�6��G+�!#e��<��
��IP(]s,� �x��$}���7}�LXo<u@;!7�g�=0�;j������5f����_�n�bȭ�b��y)��ߊ�>��K,�l_��b�x��/���'e�q�
wC_�;6{����]��V��&~Ck���D\�#W��Q ��._�i�Q?8G�������� ��ۤů����=o��5�`4l�欋`"%�<RW��,����C�b���+����������� �~�Q���������TNyl�6{��~���=�Q��Q0��=V�g��d��)M¼Z��D�j!<,2�-2i�.�u%|\��q�LX��qȘC����ߗщӌ#���ĩ�v��Ť-b.sE���� ��� �6Y+����g���*�HĠ7�&0�N�n�e��z4�dac��6a430�@GV2� (s�� Dĉ�T��ta������0	��lD�
���q�h�+2�_�M�DvX��2������MfB�BM��eЂ��[�A\ɸ�R������*��*Ũ%
��,hnP����J�}��( >�(Ƿ�aE9���Q�S��p#�+�Vs�X��υ>���4�uCM��t�QC���=gj5&�lȇ�?똹�}M��K3�+��^yb�M�{�ZP`T�l����9�G��J��0���h�1|��J8?�vӚ��A��F��� b�ʩ�8Ϯ���,s_C�L�g�T��77�O�A��=[k�N
�s&[_��0��|)�����V�W�}�z�׌��42g�V���*�����P��^�΅��j��v�C��f�'�:�AW`���?9�T��8�\h!ã�C-��>в}��UA�c�A�q�*��i�LGC�zo��HLcgvExy�[j8�	�M�V̩{u��m�J�-�Ff}3=&��m�C��{��~�h��Wb)� �Y�<�-�"oUKڅ[��b;M�Kr�"k�!�ҮV�6~6�z�O���*D�I��l�i��ոț#9���8#p�WŠ��]��'1VNn+����,��J%�A�2�t��~�̧U�hcC'rv�H??����.S �bR��?��0M[��؆�3�A��a$���(�[��� �t.�����X�ĝQ�I�\�Mq�V�{��_�FQ4^ z����C��0E���/�md���r���1������nx�I/v@%��86�N]��K���;}ηlXb��>@<��k����B�)E���M��۰��XrM}o5��B�u4ۘ�KD"�[ɵ?�I5RP���8g��<��l�|Ŭ�;��S H���7E'�2A�)�)끪���V��|xu9�t��1�
y�%="���i�)m����؀!����΁�U)��cm=3�Q�(�xiw����߷����F"�j3�E���Z4��[���W,��+��`�����ְ4iq���z60�*[�wz���p�=��T�~3� = Vh���拝���}nx�O!���i�]K9��X�:�w-=	���8Dr꽾K�r���mu9�A���t`0�K�Y�K��`��l�h���Vj^䷵շ��;�v�^�/�����hKG@��YD��iq�Lǜ�!�F��p�%�"!�F��Ж���3�ՓF�Bl'�Z|y��	N�hE���5w"��>+C�D���Ěr�w�lT@�����,gnm�y���5kI`����x��A^��!��4mmMV��mF��˥X-����lb�(�)�g杏W%p|�]��2q���Y���ﾇǱ��ctn�S��艵wj���fp[������̙S�$ �$u�������5���-�$�by�R�������i��5Ty�ڏ�����x��\�~�]3��Z5�D>��8�������n���c�Pt����t�X����-��7MD�"ǎ5����*�*F�W�D����;�	o%˄#��G*N:]����\�� ;��>�ýBq����	(���f����_a����R�[�-p�#;�v3����J���DN�'ϥ~��]��r�Р�k^�k�LQ�C�%?�e��+�{(�xGf����9?+�T����Լs��3�SS�eC�B��5m?x��=�Sތ�#��G��8%|Mפ�z.���/ՎX�:�c���hTV�`�o�V�w܁�2�
���j @����9��=�t��7�X2`�/��ָ���I�%���9���6;[��h.�;o�#��&���q�^�9#kH?���O:��@����`�}�@�3&
��O����A/�=Q�L5��Q�֢���'�����:΀-o5�>�;4Lt
��m�AtI���d5��C4�JJ5ܹ��n2w��^��EV�$�>e2��0��宂�9�~ȣ%��H��P}g]o��c�jT��r��"���e�k@�xjBqV���?@�q��+�>0YM���q��KX�=�]�L	K�L�ց	���򝝸H�r�v�5C�����IEjn*�ː���`���YA��҉�WTٕ����BnʷXn���\��=�u�#Qx��[�bJM�����%�����)H�^wNʂ����V'�wr�1�2]!�EӿC�"u���_mZnJ�K~��f�]��IU���D$�Bf?#��������d���D�C��a���I��XF��.J����ΡK ��y��4�o�ʮ;����
��5��Ȍ`d�՛ꠔ��ՖuZnO���6Ɠ�\��°`�zT,�S�Q�b���5�Y	�O��-q���:�9b�z��F�x���ܮ*���i�����y{0M�BC~��v����I� �&�Wpo IL?�2Q�W���o}��Q���z��e?i��I!�<���I�0�CV��N�H'�Gt�..���������� <���s� \f�y�My�͝�+xQ�y��_��<��x=��W`��s���/������w���((� c�����5d2���6�,��&5�K�ڹ	I�>�YG� �>�a.��a �(�{N��J����9�%�/�.1q5r�����$�(�[�ƙye����n�r��Q��q���I*l��Δ"����q�aE�Nf�=��+*��e~���QU�ߏ�aZ�_ҳ�P��7�E�=�'#kA�5VA]{i�
�;<��@,�� A	����i
��������]2�%vLC�$=�#�,�%Y6}�*�l�X>~G�ow��X����XŐ9w�oMɮgH��/�P��Ēi�8C���r:ch���\t�G/���V�Q��}*G\�����Ʈ���[5\���PJw��L�y�
��/r�3�p����^V�!�[�q��qP~]���C �-M������F�z�8Ddէv���-B�IW���~�^P���� �0�w^}�q��U�g�X��kzM2��R�B�-0��Ǔ��~��ׂ�$	��w�g���@�v�Az)�Ա�c�𿐜MZ`5�_5��T A�5?�5�`:�p�m����K��CRu(D��Дu��B��G��8����x/�w��#Ψ�L+%�D�К��eٲ|b�$舞���>�Iఐ`�^n��UF�������)�$\���ű�_�'�Rw0�D�`C_�V�j+C�R5oV�U�bϽ�>335:�韀N���ŭ6����!���_�I��9� ���krn	|G��a~���f2H���pϒ%���e�67<���aq�q�tJ*����#��h:���.u�)�f ��U��o�Юl��ucO�$ �O�n+G_<";ݹ/����v�%7뼞+�3�v������mH����]��Vnl�2�l��.��VXU�QfJ6���w@�(Qͼ�l�.WUC���u9��$E��v餷�s��gJ�߅w|#|�Nx��?����G�|�����>Q��E�<��R�.��#M8��D�mF�0����⾠�;g�J��� ��`����'�v���d�8��i8T���0���WG�= ���� ߁�=R�@�+�@��n�l?+{����Q��췮�p�W|�rA�B���})0j.Q�ߓ����2=S��~��k,��7�@������a\	;���K� h�K���(ߐ%��/�Pk�
DVvԔ?wY6*�� hu��"��Rn`W�,T��م�����~b��`@b��:%Xs-Sio��C���v������l!��[4fQp��.�5��B-����F�T��\��y����M%ϸ��{J$��w�k�3�N0I����ĠR��p�a/��D;G���J&Kp�o޼�L��n�a�=0��2
��#�=q�C�HZ<�*	:ȿh;��qae�x(�D+@'�P�켃��h�_�Z�m�C������z���8�9�5T��@.Q���n�BTeӨG�R��G�����f�-°8�i%aG���Y��=��^��W���z�<ȃ�=�*��u�p?�MU�� 
HJ೧�
PeL"�� �{@�'�x�/=~A[���� #!�0�*ԑ��
[�a�~�m�<��"��˭����Y(�@�bޥ/�l7�nq������S5���ȃ49)+D4W A9��0Ji������|��`�<ș�k{�56 ��잿֌h$v��K�$��{�;�&�N�	��W ��#�W�<����7�ʽ��(�(�X��۩�~]㢊�G�gD�p#�%��u�XK�O=Fa���%#���c�����mpmp[?݄ �fj�HaghUG6���^O�{	,[�.+ccU-��$����Uj�N�A+$�Q�b�
��3���.�ÅKtb����Y7:$>�SE�vXi��|�wIDʰv�]�X������[|m<��BǀSI�r����,y�K�RE�?��]>�t�8�".���M
h��)qh����?���]lN�qŞɄ��%j󇑏�:9�Q���\�#�#��
�	9��Z�"�
������ZM�oU쏏��I��J����G�zWo)�� �N|�|s,���RZ���v��}�ա�O�SmTi���_��Z��J��2�tS3!��a#�X��ʠ?�4�N}+��F>Vo,�M��;>WΕ�����~�"#�t�S��_��1\��(�^_ۥ���l�����pi��7,,z�f� �e����龞'�W�nʳ�}�D��y	��^MC�U{������q�e���;'���l&S*��vqE�Α�6�di��i^OR �6*ٻ7�cO��x�o�m/_o�zoݥ�F-i�v�|Z:��5
��{���3���Ss�˅����rQ��)> S��1�M ��xW������TC��I�c�V����_����-�m҃F��b��-�B�o��_� �'��>��鑟�uVݛ�Փ�v�_{���-4VYpp�`MP(S�a�ʙ.Yɡ�.�@i�;w��u��-����v�����<0mp$7黮8���)��0",�wc^`���r�7s=^�\�\Q�e�&�u�}8�&�	ѹ�>����lT��
�Z�RRw(3J� rI���Q)Q3#�TV̋_��kj��9���h{s�7u��E����#T��y2Cp�^qb�����t�U�E(�b��r.��:��I�x67?�{�}����<ԍ��wP�s{��׆�^�x�I.X֪���SR^=JjT~_e(�
�4��+�?ԡB�E��"���(ݼ���B]�ৢ���)�>^7�I��_�+�+$�>5�6gZ��+�Z|�%�ũ#��0=j퍝왝����t_�:MB��Az��$-��jz���Մ5�D��4S����!�Z'6A�����؁���:vMn����п��袐��ҿP#��X|�w�dB	XR #��R4X������߄ltjY��5B�k!�FbB�xE�Z�Z��}��5�;t)�mo*$���&���NhZ�ɺ����=B��ݍ�Dǆn��l��"ă �L#7"a_���U�-��-H�7��(|�UBo��uM=�BR����D"��Z����Z~�1���ͼd�K����o��Z�m>��G!X��/�S��k��5��Q�6"R��A�t�����d�E8�F咫��=��?p�@��K����4!���a�N���B�B�<Fq�)���AZ���@�b��tը�2������t|�\8��L"Q2�I-�(�,�[	e���y��:m�k�䗛��g��8���iwV�ɿ��r LF�(߹K96Q���7�B��op������5�������Ƴ!a[�#�?�\�n;	?u�v�+U ݼ���f&`�1� ��c���@k��-�4�.�O"�<_ U�W�+�C�,�����{2*t���HA6��=|i��fm��9�-*"��'�79�t$#���S����d칦���\L�W����E��PR��P��CMXv��[ǧ�W�A��U��0�L銰A��#И�\ը�Z�ƭ��*.�܋`%x�o#����(6�V^��_(�&�4n
����'�Q��gE-���a�����17 RE-x�UV3tnVL2}{����-R�z1�y��cGW�ۘF�|Կ��>�#V餗jbF��?"wU.��``�wIH�ޤ
ŜKnVqmO4��@�3��=��{&������w1H�P����!Ҫ6���e���.�D�C�u����C���s�sR�I� �B����oݗ��ݺ<�^��ƴѣ�d��gѫ��!��K.,6ΛM���mS��Qs��C,"�.���z��W�n?˩Ñ���.3Y��#΍�Pp0�$��p��n��շ������ߑ�{�&�����A���,���%��%_�T��|ח:8$F�`��>��R�;4�^�~W�����4��x�W"Q�ͣ?5�W&����ӏ,�)��% d�R�������������-���,���q9�]5��s�W�0�}#��Xac�6��x!�����Z�
5]-ג�������a�j#�3��}��é��=�+df+s\J�����Ե�F��8��丣چ��Yf�qyg7��F��Pf�+�1�9���,�Xx�)ݩ�(w��D��0^��)���ҝ���W�t�#$H�&�U֦����2@j+��Ɇ�H�f��)d��nH8c��~fbH;�c��۱��5x�ku����X �n��V'��d��Z���u������G�{�[�4�L`#<�`B�^�_cgc�bҰGbV#��}u���B�{`7ڵ�C-IX&�'	5���p��˃��u���g������.b0%��gZ(7���D�P6���D> �i�궿W&��/!IZB��Щ_Ug!��0h�i�[���3���������1�f���2�C[�JX�%-U�� $��&���AX[H�ppť�0������eU"Rb�*K�R��6G��ں:�D�]Hm>�j�E��=�x
\�s�)�C�&�!=:!�ߴ��.m1 �_8�,�:q]��|�Qދ�pIڵ7��cj~O���"�B�F��mf�W�֓nje�/^˽?"N�������$��C�����*�Ə���UD��uݰ��#s�}q�lU#?B
�������<�e9�/�E��>P��o2i�^��	��܏�5�����Xh^��t���dk,%,�Ād�����BKj[t��~���ᏽ��}5��YX.�в��Kxn�;�)Uz���0�)Kę�_^���q��#�"@ۿ���jp#5S�@�:��^X<є쑕c[,������)^
���6�-��~	�wQ4t�~�]�o2
����%�bιKl�:�:?�;�X�i�f����9��(0/�q�u/�.�UCۑ�5�dbKf����7�K0ZQU���S8���Q@�ocuT_�����v=��x�Y4��xM�D��+}7w������g4Ka����	�e,ʯ��o��c� �$��Y"M���]�G[3�*�ty��j��-�k�;*+d3����=�ZH�!�QV�Soh���6����]]��;9��O���A^&di37j"���&ʆ��%�+��u�XӾҽ)��P���ٙo�̔�Jɑ��1�2�5|E0��E���#r��_@�ctwg8��#:l�V��s��,��X���׏3��	�nNWL�LϜin5M�Z�$ ��/"�mO�ͭ@�2*�S�!� Yua�s�� ֿ>�̻g&@�>�%��t���F´��Q�R;����_�7p���7�
�Aц*���%�f�`k=��β�����A'a8�{u�����:Jđ(s�W��=�G0龞�o5��f�}�<wj4N�w�s�Pğ5����Q�ϫ�؃IK���1�n}fe�)u-"�U:�LVҽ�?���n�D���sD�+_�?�����+��!�4�i/��r���u��YP�fMS�Y�������co2��[֢+�Q{Uv2��C�L�dA��;����z�4`�H{{ֈ���CF��8�:}��'�A~��x�P�Gf7����h~�U� OC��h��w�<�`Mf�g~�#�;OzI�;��
�5�����pk�0��A�1�7W�Bla��-2L���J���1^�SQ�B�q���������sp*��M�M��6���˷>އ�.]
ݐ���0�:�L�	���$bF��CLYPn]fYWD�{��#wQy���y��`�P|ޡEʦhJ(U��P9��$@�m��.NQ��Z%�iŅ�dZy�y�C�@N^(�)��4T��7a�� ����ǳ��&��
3���&N9Y+�����p"��?�TRH�R��tL의��+'y1��������q�2��Z���g@�Beq:�]��!��-��i6mt����w� �b����`��^���j���;dY��Z����l�ޚ��q=��G*�f���F��6��wٚ�%��%�ݒ�4�@Pq�2F�?H��k(��LW����-j��	Xݤ���I�9d��|�W�e����\�|�سI~�m��՗Kֵ 1 $g��q�dZ �������aL8�,Dy����5�f�e�^�?""Ǚ�<@�,�A�-0�eA�psy��4=AZ��Ʌ+�-�W�~0�� R[����:b����g!�������u?Ԯ��nxļ�W\��O�<r40Q9�����X����l&OiK���k�� 2x�~�����b�x7+]�\�˙YB��3l�1/ĝ.N�-dTvg�$7�����XL��P&(Z��\ō����*��}\��7ҺY���Ow��^���Qt��� �2*���y�%���m��JO��)���a���qQC����ʨ�\�\�)-OM��y��7K�O�\�7����*����ڹ�����	�x}��MϮ��.4b����c��
�bQ���I/p8hE��*]cd98OcԼ�T�0;����X�b���z�DY8(;�?���6�� ǉ��"r� *5z��,u��\�ք���B���,�-�1O׌�~���h�HiQ������.�ee8p�4g�}`�`�X~�8���iجi��F�k��v�(�`���1�f6GMF�����N�"�&�_>���Ju�.� �N���E��A���h��g7PN�憊�&(ޠ�l��� ]QP����
��2"���#���I��� �[�/#�M����U�Z�^G9Y��#�_>V#����<�n�ܘp�OT��ǎì���F������\�\�c�����l�?s*s��v�P�3mU߷B^)'�Lim���2�D>��8�R�	�֏���?&?�2�Sz����R[�e��kH$�ݩ���9�}]����`@4.p��6�_�GW����K�C	���A��n�9|A��$%��U|2/���DQ�N�7����-�����WKΚ��-�l� [��z�o�������QD���+��h�v<Ype�+�������ޫ��J����GS����k�x�����װ� ��H��Z�)_7n�$�ǍĿ0��dh�'�;QD�k5���O��nF��g�Tp���D>&4��eN�pS�.�s.��E��u��-�ƌ�^糛���_y�,�$��1O���Ni|r��[
�+W6l��O��l�M9v7�P�B���,/'뜶�IUm�vQ?d3`��)�&~%��?Hyx�/����G݇��}����Mr,���:���|�g�ޏR���@(�]�x�]Z%R��{�WCPȢ�y���L+��U�E�M����^��
��!�tq/<���b�Y����x�}��ׯS�������fͤލp��X ���hs��GNE�.eY�0Ƥ�$�/qŵxJp�kR�N' ��*�k���X�T� �I�S�6G�ƽp��t���Cf\(�?m"�K����]�B���r����_2;E�%\s� ��#�O�-~g����[I��a�r��K�F�gXڨ��7�~I��}Z�ゟ�)pN>���}�E,��f����4����%�(�U���*P�N���{���R�<	"{<��s��ʔ�7���'_�Ҵs\*�I����ߑsh(0� +Mkl�k}������a$3���;е8i�;���2�c{� ����2�ڭ3�e�H���;z:4�Ie
$��N�|&!�� ��3i&�����_>�(".rLҀ��x��=��G�>�D:�v�7Z�>X���#�Ly��(q��td���A�>n;�<k?S����ת�*.!T����2ra��s����,R�B&^u�o�>���Kˌ�	p�v�jAMJ�(���#��ۘne���a��&�~_��?��� Y���wR������JF�ӟ�_L���T4�����E=��2yYG�B�gGLJ�"(|��Yv�$���TB��Sߘ��	�"9�˃*A�ԧn$^� �葁_lm��]���Wn�#3cE]��E^��\BDs0jR>��]���IF�Z)��XM-�%a�\]����JS�#XS�7��	3�H����-�p��ֱ��ݳ	V Z���5�?�d�A�Zw$q˘z"��g���8
$E���Y����� -�<�Z�\s_P�� �3��Q����&+t��.��G_3�1aBX�{�����D�%w�}�x�@�2�/m�p��]B���4ń��[-���iF-8w�1%I��T�X�_b�D�߭��w~fh��:K���>i�
�~�6�cJ4ؤ�ó�I�qJ򱲢���*�M���N���+�j���!��[&�TNR�%�t��II��y�#u3Ń_~�m��1v�D��f�߭H!�)���(<�o�NE�@a��a�f���?F��o�yE:!s��|z�pt9��w���SL8��ę�m2k�oCu��m#|�1�Φ��4HD���{�V�U��iH� �@?��[`Ac��M�#��:ﯓ�W_J�[4u�!&Sf�9�n;:��Ŷ���D�c��~� �(�OM-�u�#K��a�a�킮'h�w"~��ݯ�,��>G�B���1x�2g�R�ױ����:�E~@��HH�ⶉ{ݺ�X�r����!*�_�k��|?rc�"�Z���>BV�2���#�m������3�_	���D
VV�*-�h��A2�f��bZ7��H���J���v9��8MK*��Y����W�͋�G����l�]�y�{
�}��A��n�ZGgU��H��,u�ȹ����P�d?�v�o]	si7}Qw��`�N�5"�q�!
]'gɎ�[mG��2)#�#��d���&��,�s�}���y�`�o�j���b&�.���H�P1U�.�p��7��Gg!n����_��3HEcÜ�vi��約��ӂ���$8��?j�����(���<YӉ�g`	�C�?�R���kq��/�%�:�r�+K76|��V�x�,��j���zR�Xp����Ֆ"���p��ޠGٟh�)c��g�p3�m�P��Z�4��Rq���;\�
���1�u6(�uط̿ם���De�Do0H��\*C��.��Y����٪���G8����!����Ye3�����2.�Q�o�Α|�|´����~���I���d���zK����b�����v$n�b��@3��|V�\����L՟������Z����`*��)r��e>�:����g��v|����j��0���R���JY	������?�$αεd�fl�AxӀ%߼��*���{�pAC�� J.��k
R��!�;bG\�h��b�Nc�@JF���~��@�5Z��-�&�f/���B������OP��,i�a��#J��P�ձ��y�H��g�XD�3)����l�R�a�v�e*�g}���0�TG��$�4 W��)9ގ���1A4�E��;�HY�����U�ˎ���H󵏓�]�H���b�ƫY���B�֑js�3� �J� ��]08���^̼������?K�A�=�һ>,��[>���EV�_(1` 3��,_��	�l�����
�������;�1�"�$KE�e�v�]E�R�a.�tea�A԰�x�s�&: ep�>�h 
aoر�͛�ޜJ�����fܿ����,�[��%?Rמ�c����B�I��:+�]�KP�J�ƃ��>H�5?H�p��dM�r1����r��|��@�3�7�r���&�q�ы.ti�x��o�B��g*�TL�u��0J��E \0���\2��mT�Sۿ�L?��w��� �����a,��Z`5`����E4''�=���'�
�/%2����N_J�OS� �o{֥/��ωO|��O�2�I�J@�H�VR�5��0Қ��;�	T�K�<3�Ⱥ�׃�T�Xo��l8�Q
K���o~FB��S�;�
A�LS�\AF�|���a�#JX�r��sJY덚dDB�Q�o;�$�jB�-�W������-�=�^�'�,�|���tK��#j4��ӻ}��kL�Ha��W�a�q.T��n�&"�U�;-@����<c��m��G����d���1m���*�F�[�G���#����qQx>0:G���-��zR�t�b��'�� �FB�K�F��X6�9�C������q$��s@E)�x����W�XŎbL?8���|��2��sάv�[a�0CS?M�O��C�f^��ra���?�J��&�OȻ��I5k��;�%�G����l�(%�ޖA��(Wνv�V��F7v��h|�@����Z�Up��<+x������J��c�?&��'7ω�ˢ(�I���������q�ܻ:�&sb���������S�.�k�i�7��9�eV�;�0� c�����Uo����Ih�'	�g�D���9ܗ�!r(��L���3x�ٲʬ�sw[����vCl�dD���M�@��� h�w�	(ȫ#U�4.m#e����DF*��c���
�h.l{ov��>��V�&�v���M:}��Եk�S�m��zlj�����T:�i&\|���������wC�cp#/ǵi@q�d_���Q^��_6��dB���T�}Y�CKa�:����J��%x���7��x 奯w��T�����$��~?���Hn|3_9&3*�x%z-����Uة�A������&��ǶǺ��glk�2nPS���,~&���A������Fol����E�H��*������i��qZ��`ӡ�4y|QB6���u�N�:-[��շ��{�daSZ��>�%Y��p��p�-�U��E�9s��Gէ�E���2M�|t�p�s}�.�������۴�)���r�5<v=�#����
ϟ��q���;yp�����Ƃ��K�Q�ī�2�x��ڃ��m�+?���r���N�bsPy�iv�*_�w��CU^���s�w8g�]��֩���=-xO�6�і�H��Ɋ���n�Q��L�G0k�+�>�ݣ��S Y
}[�dx�Q��7�:zb�*�B��wY���A0��C�bf�P�	XBET���]ʦ-�
a�C�k�����Jolis����\��Ò]���N�YsDօ����dU�:����x0�*Ñ���;y����ά�ۊ�E���F~cNe�MF���p�2B����/\�}���A��a�׷��?��Y�=+�Z�GY]��jt�O'�*6	�u9A�v��zw��eo�7,�e�ؑ˴�D�r�陪`U ��)	к�Q��s��c�W���l�;���?l����JT(�U��p�o�Y��O��N�[-#ᕩA1���)�����p)&,}��Ʋ��Xus򯺏IO*נG�=��$�s.�H�웩�F����HS���6{�`����Y߇�E�MH�VT�\�C%�w�5w@�|@|��E��b�����Z�jvwC3�S�=?0*�^	g3��؃�%��WQ%&[��=���*)�]8]-�~�ܚ՝H�_aY����^ԏ�yt���8v��[�6;��7�N)���&S�:Oq��:2�m��FCB���ly�פd�5j�u����b�O^s����cu�4]xf��	���WE��X���b�x\��Er� ��*�
��BJM?�7T�LSL'`�ډj�J���ƺ�5(%��IK�{㌷��`��a���р;���W�?��׭�U�C�}�%�s�G}���KS�-����+���C"�]BiCh�=@\�$�_��oV[#����M8�h���Hܵ���������KO�V!Ga�h��E'��2�r80 �5��\g����V�+�Z�=�=�Os���w���B�5�?��������6�O���@�!V�����%�&z	B����nHvd���GS �6��kq��&�����I�g7� p��Nq��S���}\�k8T�T�s�:�pT&�0��^"m��j\g,�Q��0\(�/�	!�e�*��wk���Iª+3r��2F7��?�6�!����#uL��`����X�|p�	��Rl����!��Nw��x���2P��RC1�)*�EH�G~��@Gؐ���e�K?N|\��o�~b��z)��fʹ3.<d3�t��-���V�*�Y���	�Q���{ʣ�N�R�E ?�8ڣ��RB�B3�5<�����m(/��#��"�^F[S{9dp��"�����p�<�eC'ڑaǣ���G�'��H(a������^V��EL2�ȡ!�Ob���(�A�Ȯ�#����פ��ї���q��ඁtg��q���j�%������6�	��7gDk�m�Ew�$���a&H����� �	zcS?K5�>�b�N�t0i��������V^߯�� ��1�z���w�S\�E�e�H�'/&�&e�]38窉�^��p�r_&�
���lD��W
�`���������S�I=�B�C���\RH�P ��զ\yZ�Q��L�SU��mI��aj�PƯ�� �˕ն�du�d����٪I	#�m���no�]��NvNd�x[���nlu
�k̉ ?����X�ym�`5�	�L����|�zJ8-�.��-:�Q/@��J\�}�'�tk)�/DWP�y<w4Y��h��j����B��@Ѿ�y@H^�x<�h6�<	Q�Ĺ$�*WN�����B�|cd�}�J��`�sy����p�H�VR�6�]G�i���nl<p�|���'�4��֊�QJ�e>�^�ސ�ӊqX�C�)]�`i�7����@��1���/p�%�)!�.��Cpi���P�=�0&;�/��䝩�O���qꯐ�I�$�0u��:�t/��|K��e<h�9i[E_�[n<[[y���)����Jt��?�tc���g	.��eA餌�n4��=���؋�o�>��0��Ӫӡ�B����ܖ��i�WdJ�ĩg�VG�;���b�,��/"{�R�c�c�4A�K)��8���,��W�a�c�n�$�.&\�)�2�����9�Y���}f7ԍ"�o�c���;wkH:؛�-��=��\13QDk�Ԛ�/]�l��i���d[(����ɡ�#���\��ą�c�?�~#�ⷔ�����I��͝���#�U�@��uXXh��M����7�
4q�_��?���/;����T7���,Xc�x=�3fI�&ZO�蔯D����:
S18�` L�ϲ3`��Ϟ�ey+��A	}Ç��<7-�Ǹɟ)����I�Ҟ��4U