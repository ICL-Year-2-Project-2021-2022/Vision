��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�
TB�(+�
mQCJXA@�A���k��h�U>QF�q���Э��f��y���W�k�2�e8C��:���lO�*�·����[�f;(q�i9�Ҙv�,v{�@�gw��<vT��əI�2�,6�2��I�n~�v!�y�����O,�|L���D��L)�$�ݪ�yy�Z����Yj��h$gQ����8�Pe0�!��A!P���_�Q�T�3^���'PXeՍ� ��SO�k}ѥ��>���;��^_�-Fr���#GR"z~m]�*�$>x*�a�4-�D�����[�ٰ�7�&p��,��ro�ޯ@A��_�B1��:��=�&�c��z����F_�1�(�l�<�L�H$z@�b�=į��)��8;&�k'U(X�%�>� %�22B�+���j��7ܯỡAs���irؖZ2Ӫ�\�o�PMj5�t�����u К��Ɵ��?f��Om�=PQ�g
�[��f������$`�ř����,��6=��zRl������x���6�x�}�s�)�LElE���}�*���f����P�}@+���$Z���y��H���o�9���Q�?����֚1����s|!��Q�����o|Sgcs��̂�=���G�
���-PiE��.�5G�P�đ��>.�yçZ��ߓ/���_�"I�>���'�΄����%�x!��ڵ�}m��0�4y]�H5V����Z��S\zj�$>�+����U��Q�jG��Y^Z�R�K�4!