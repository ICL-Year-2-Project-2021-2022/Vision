��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P3K��$�?~������\͡��dk�⍥xm3T��8�׬����:@Ӻ�n~��6�*ݚ������a4�**�1'wO���?�N38W�'�T�u/���~Wpm�ك>p��Ѫ�=��+���Db�$�|�^h� ��U�R��b�����%�P�gJf�%��kza��>�̴���͊��g^�p��J	Ki[ڈ��:.gE���SNw{d��S=Rى����;0��N��t�բ3|�LB���`�F>%�����4[ro�3��+���Ƴ`CQ�����NGA�,�I��11�5QWӟ"��ʠ3\�J�*N�q���k��u��ӱ-΀����w��q�˸(­S��9pZ���h&%7�����8\&*�%�]>��?)l���5��o���]LWw��ڿ�a��܌�Z��ټ�8��7��ZjM�;�*�B�� PJIW��n�Y����r�4^��Lq�]U!�`�5|9�U��C`�@�j\ww,�j���Cח!�2��w���:|H�/��0�8�����3��R�e����`�z'���#X3�q~o�㱍z��{��G2��[�������[�*�'%Z�\�t�����������jӍ}z�w�2hv��h����[��br!(��#ѳs؜��#FM�_m���y��^~ԇ*�s���M,x�b�+m�ޤ��xտ��G��\�:/����7����nU��A&�Ml��E�DJԆ�y!�J��ym0��fdmxV��K`�G�C���c}���c�ck�#Ƞ�܍�>η+��U�X/+L!�]26E�g�S5��������\v���i¯�Q��V��r92;a"K�)%�r�9)��B��s���%�i�Kj���W>��1Qe�c�*�Y�2�}��uP~���"�_v��թ��`4T�W9�u�ߺ��34e�a�{��7�ɥ�<��~<�n׀���$~N룫��-��_�=rG����7�16�D�����7i�&��w�ec��=\��2�O(�T2��(�9����BOE��[�����lɃ׵9-���#tݠ����6.�����Z2��]
�p��FFi���ت?#�F[%�x�"xz cd����L�B�M
{�@8�������X/	�ލ�Aa�T+��ok<�:��B�f�c���B����b�޻�0G�$�Oߩ��AZY�����|���#,�Y�S�=�!�jp��]��V�a�g�"$ښ�7���z~���C��·D[3�o oA�Y��D�0(<4ޔ�g���'y=�����m�S��x��2ӱ�'�C��z��sVp�aa~�D�p��3�@��'�ɴ6����������_��K��( ��쟠T�덛/�>�O���w�ҹ�j�*�b��S"�w
]�~���Z������o-zӾ�\0�� ߣ����4�����c�F�����	L��}�U�.�G��"!0�6�P�<�B hG����2\��]��/��"�"4�}
1�(w�z��x��.�߱H�鞺��dH��W���T��7c7V�H��B[�U�� "���+�Ð�����R:��F'�Ÿ?��%������j�j����Y ���-G��{�/ww8c&c���c��Jλz����G��-��y0RCP�����\J���@G�R�b������$��k�gN����R����ޔHt�䆱����zRi�"���K�+i|����PW�cI���`�W�ѓ����!���z��&���沎V]�� �-"k3���W�k���������6$N
��t��F2562�E#��]*��o�3�E�ױ�D��T��kĩ2i��A[�9�ךa[S� �hw����_@�ya]R��[���"��������^�(BJ(2-���e��N�� RHLs�l��G�%��5B�
�����V0/?�%i(�4*A�N�oQjaВ�>D��4q�Jh����?ڞ�C���;�RJ��HcWmGЂ��aC�.�[f�'��\P�ONal����(�6�Փ�Lf>
�L�Ɔ�&�{����y�ic�F�\���O��Կ�VTt @Ď��,>sM[>}���Qَ:��Bņ�t��������G��O��_�0�l~!���L�
^QaD���L�
��{��Gj����gQ+q/E���D$�=���4"��'{!��ʪ�AT5�bD?��n�+ԍ��^��^]jX�8�p��Բ�ɍg^�<��ga���Fi�Clb��YO����35���� �M��#�$�:ZF�ͼ����񈹇%Ԍ�;��5$�c�$�(�j��́�B�ٺBC��gc_�o6m��>����������
�_�h4�(z��(�B`�ۍ��"�_�$�]���i���fꜮ+�W�����/)[���mf!�1�-F�ّ���I� ����*Ϊ��yAm���q��*�m����#���{c�21����U��t&z6��s�/z7b%qD�B�+՜h��໠m��*������<4v��J�K8�^5�������R�l��>r���~$�,o\�I���{袭��� M���!�+7�b}�Q^�r4,1p�vHL���Ø�=~9)�~�+�H=�3r(i���xάEҹ�/Lg��a9G �(na�(���PG�LBER��]�Z��P��^����-8�C4/p��x�qb�y�%��{��c[��m�/m�]�����'a9{vlh��-��+_�_��1��<!�}(��w?@'#��D	X/�HE4b�$�l��X����{��v5o2u�78��~�ޠm0�?���ŲX�J)�t��2�m�ӈ�,1�ı��D �8�}xP2�KxWBg��m,"��T��4x�>�/}*Z�iN�,����D��OY��H�`(�&?G���3X~�cl�$��u\�ǻu`�����F�Nk�/���.�^���mX@}!���nuk�u��-*�.��.5L�O� ��y�y7�*7��[k�����*Нq��	'UR��[CӉMot�N;�z�+�D�7�݋V���#�si�\[L��Ꙣ	v{�U����1K�;�O���pv޿�T��b°'��+��a%y>��ȳn)�W�����@�`�VA ����v�9o�nK��T�z�(y�'V��5wjuǹ�B%D����qx����N
�$1�ɰo24�"���Fҿ�J�w|�뎐R3�H�"�����s��ȍX�/p����$��eѳ����X-V�"ި�( �����hW��)"_�J'Iwn-��,|:&�?����iO\fN-�����sm���𽌄|s�����L*4rh��?֫-$�_��%?��ٶ0&_bkw}K���Of�p��q�W���|`��񮆓��%���p�����ͬ��fY��.��:�.�#o�s�����;����
v �^�EuK�Gؿ�"�c�ǾR�"�d^cY��Z���#rZ�0T��k�3��q�����d��t"s2�$�W���D%��D5c_��$��|x�׶�t����a���^��Jĉ"1D�X�zt��+�OB(�m/O�@�N��h�@l��!d��x��1gy��J��)M=s*�5���Ɖ.�e�r�ӕ���[D�\A���qб��@.�Z�,'$���f?ٳ�h��Ɔ���pP��Q"���zYa')���:��L��h)�,��>��'�m�,��+�h@�1 7���e�w�ܠ�O�]�K?̀�cs�d��[�5�;E��Q���('.G�3]}�ɷ{N^����)Id���c�4�l��U@ڻ"ۉ�)�_W~byd�������(Z����?�6�/eF�D�ˍ��u��Q�:+qz)���š��]����6 R �dF��P����lh�PF\�j�24�B�}Oex��\/��=��J�[
}-�R����*�����Wa:
�:xTȁ%a���"����pOš\��:M�����N�e7n6�
�A`m��2�9���|xd���>T&�$&�O��e�2���UEe튭Nt�`�8���y..'��}Xc@}�M�#�mLa�C4�sL�'�'�V����~���K�Q�-�\�g�����y�Zh|���.���e�F�ncb�q�3�%4΂�>�݂�^��m'Y��}��?d���\����{�.�d�~��E�PIR�A��K��o:)�j�;o���'}�$T^���Ē$NT}-��.nUq,;W<���B�'�TYm	$e�3�>b����4�o�Yv'u$��'����и�"�bۼ[!��&`�+a��c��;JmIj��u�<�Qm���xl�����'����	��!mN�P-&�X@�K�qΦ�v�+-�|	�+�4�q����Q1r-d��0=�f;�j�`�M�����B��~����t�Ɠ2�$�YPC�2��F�X2�K��@Z_�\��ub�m�Յ�˷B��E~�o����]z���0	Bz)�$U���l恨 �@�2���خN=�֛"yY�zO�IÄ���
� p��s�ms�&6���}g;�"���e&�wƿF���䐉��!N�K6*��0:��$ l�c���gvN}��d7�����f�SqЍ��� �����g�Q��\*�,��#�,W�XzAR{�O����
31�P���,ٺ_�-6�$?��t0՟��0]�L�Z��S�i]6�)2:�6Gw�i_o��!��4E_$l�]P��Ӽ��'q(�C������@R:qA+����EK���/�����A�]Wb�;V�__���x�	Э5���q_���|�O~����Ѯ�J�%��b}��)lF�s���9`v�HȪú�����4��2�ci�����'����U���lv0�����8|�vQ,G9��xH���}^X��j���Q�7��u5�{��a��ޙ� ЊQ��A��E��-��L��Ә2�O(M���Շ���j.v	���60��Uf@K�KK�(V����Χs�G���6�L��#_��@� �ÑO�5�'|��Bm��ch��zX0�0?�`;�����wshz����_���:��'�ݷ����i=�.T�/�R�Q��c})��&̺�UJ�vQ:�0����CpՎ�S�\�x!���G��W"j�ЉE/4$�	f���4��E�O��ݕl�4�,��}0[�����*u��*{�w�$�Ȧ�i��^���m��RC4�C��̄I|�7a��y��|KS�g�35���݇M)g1&��H6 x��3{���M�-mK*�#f2��9��_5�س�rb-?>���T\?	���{C�kg��c��Rex��:Ħ�Sd�d�I�1�T$���@8��1���_K8�ȨQ�5�o�b�<x��)��6���B������x�SÔ`"�F���=���7~�Â[T�G1 ��+�N��|��v� ��eJ�`�z7G��+ސ�6`"��1υn�h�@��7#�T�Ue�� ��rjDZf���0N�fPn��,m�I�n�k%��m�Q��0H�s��EBy1-�E�.��陴{��N�G��&?��J��s��/)DA+�y���'c}O�ra�L��|��-?z���׆�F�mx��	�C�K$�A�b�~y�z�B���G~OUA��8*鱝*�w 1����̈́�;�Q�<����&�#�4���o�VIq��������h�Z���i$O<�ɻ�S!x&��eۉ܏����DWY�M'�i�G�����K���د�L�|��<c�w���0�"��0hW"������|�Ӽ�+9�ǂ��݄u~G�㴮�Ö}�|�c�Y.'$eg�RE�qH�������H�0�$aA��L�G��)�z��C'5��wrBR��j2��lF��'@�)4=�@�w�%ǈh�y~�gBM�����f���(P�)�1��fo�!z67�zǙ�ȭ�S�f�K7�a��6S�F�X[�<!Y�` �w��:��ٸŽt(>~��1J��G�x65)z#�"1QlMv�N����8��U�H���p�j����)*��I�c����^��\W�t	&�m�7Oz�y�q��*�qn#[p$���LAd�b���/+Y�	,���Qc��N+���q���ځ�����2�Z;�	}6�m*R�5�_�ҭd!I�T�כf�>(�Q8A� 	��JB��R'3�����q�~�d���(r���I�#�j��,	�V��f��ʷ{{so`vH��2�ӊ�9�4�����5�r�Y �����iՒ���_�G�v(�U�G{� Ii���Dl������s�RL_�Ԝ^�	�k�@*�R�T�[_�ԘI)�H���Ԫ�"%��& ���E}y�C�k������P�����������~�
��$�M0�3CK&o�L6�N��ޣ"9�jpG�H����6���G�K���%���#e[�� ��7!�U�����l.�j�C2�����Epm��E	���?Vm�Vu�@��04�q�N`SAel-G=�f���^����G/���^O���a7��7��Y�n(&�OSRcQ��򷜬 �d݃L��-k�o�e�a�����O�b��sl�,�wV�:Rt�C��G��0���<�6=�
���5ϼ���|��{D+_l�PNP>���U�T�.��rP(�O�o-(mt���o*r+Ɩa&-w�
f����XHl{`�Fˬz�0�.:�p�Įq=�b�y���g�jӉ�޷�O=P��z,fc����O��1�RX�ֵhU�^Jd�0lR�r<h��X��p[��3��yM�'A�9��
m q��pH{�}�9$�V��:���-p�mr��N��ߒ�1d`��n�T�P/䊽d��S�ҿ27m�]"��Sc���į4��r��ɇ?À��ف�2G(lx�@�37�$�^O^�>��b=������6��d�l0+f���g����`V���M�آ!�9���&D�0��&J(Zo����o����!jw^:2s�o�Rb$��=vG/ %K�ű�]k�k04>�4flVL�
gh�ƨ����Y�w�H|��� Ș� �
�?��5�4Sg8G����2��sWV��LME_?�۫���@4<�F�q
\0으�)n��\��^������{��<�Ʋ�Q��0,��[ʓ��j] ����[o4��bF��`���*TKL��� C�E�Ɇ��ʷ�������BB�g�P]; ^D�%*�֤����H{#db'9b�MDk8b}��a��'�ԫ�	CNE�̫
�]����cGF{����l�|ж�2�"q<���ݡC0�F�]*e�Tz�lI2�������kH6�h���o��D{���M���#�
Ed�3}�4t�]�	AʐW�Ӎ��m{e!�u��ƣ�NDpn�(>���hhGǎO�Vq��w������,�����e���m�i��^w3焭����aN���f�K�z�e�ye5ú
Wˏ��r22Uv������12��aO4tO n^�O{ga��c�����l��X�]RJb�rz1«^0�9�t��:�%K,���Y��w��4Wv:՟6#�����5�"ƅ��+���h�+@o�Q�-в�"L/����k�7�D	��A����d�3�]���9?�������t%�'&�� ��������ok_Θ��0r�tXB�^�)QZK�I:�y��ػ�0lh��"f5 {P��>�y�	 �q�#���;�ΰ�$�W��25���7O_�,����
��\����Tq�ڐ;�~�a(�k��31ʮG�R�dſԜC]j�HFLG
Sd�b��E��[�B�rHJ�l(x�6���^���z�9����(��x�KLz�z�A�Ʃ�<x���{z��|;9C�S�~ni������;� )
�#���'0ì����ص��u�%��*��O�A�gn0����g�(Wo<c[o,B��~���G��Z���~�@ٙ:�Ɩ�tJ�U���Vd"���C�>���W�<�=@M&�-����I�5�A��1}-���ˊ�s�L�/���gLM%G��砵"�Z���2N��Ծ�#^[��G��K��M!�ph]:V��M�o�_M�n8r���mb8���BKf�;	/I]�op�TT+��������WKT�+u��.����{�f�SL�(uD�z�%/���)��x3��2�m��u�YV���X���H��j��׊4`��8G��i/�Y�;A�$9��0�[�4U���x1�[5n7f�	kU� RbRO5XxCM���;f��JdM�!�ļ�亓�i�3�*����q��&zg�i�(�9J� {s$�"��_��O|�c[�奸+����@�M`��p篆G�+yiw�x˷�o)�����u5�<�A(^L2`ݷv�f����fڮ�<�{��\��p�kXQ�0�H&�;��^=�!���,U x�5���Lԙ�ڡ��󰇍�ƴ��d{`>��3j�<��	a��w<f�`q��N�9��\�!z����N�^)n
���Zٽ�l���ӝ{��gu��  et`g�P���xBN	��5oz���Q���L��u̓��ԉLm��悇�ᨚ�+@�>���dty�K�03}�=����g����>��&�`PGVN�J��K3Ol+w^���d��6Z�Z�Wn�_��"D{�T^H)rɢ�V0�Vp"����������q]{���$!����o����LX%\�@����uG�#Aw9@۠��� ��S�i��d�o<�r}�P����I��*1\�k\�,w����_9a���s�1��u�eY�z�(�&WO'O�h���Sdݸ�_=��Gg�Q�sT����ðmx����"Y l@�P�s��N�ΐ��y�����(w�<A��!=��A�G��)V�p�Ȧ\ak��ҕw�9�	L0�~��L]RE��2�R�̢%Ղ��ėm�Nf��T1@q����W�����/i�ލj�)/<u��:y�(4'L�G&?�8") �r�,�7=��LHӋ�_��҃�V�GW��ͻ!���Q�����tQ������n��˕r��Y�����{���:U�^j}Όڬ@����(0`�+9���`K�
d�Q1��Ǒ�����h뤳m�'9u�H+�u^�K5�!�1���b�+u�6zB�?��0�!!,�F�"6��
�ξ5�(˳�~����l`߿^��:Դ�#<��hrue��xK��Y��tq�n<���\��� �JK`fH�H&'���%R����.{^p�xHR>}BL�4��;��d��VU+�2��9�|��ML	����`M*{��0�둽!x�s׈n�����(��z��/�1�;�,{{��8�j h��>#ԃ��Ed��D�P�C�F�X�8�3�zޓLT�qnD-�-����CzGn��`��|���_K����r��ǹ}u,�@j��6Y		��s���;	RE˚��y��G�шpL�j.j����T�K3�sk��70��n��M����z8�IϹYeXڱ���GF��$Ԯ'}٪l�$�8�S݃�5���נ��Y�z���|5�&%B�f(˦�S�;� �/��x�/�5%�F��	FQק�X�#'_R��|�E��g�S�K*][ư�|1&a¸p1a׭�S��5��x���`Tӂߏ-gm��a+Ȑ6I�_��/7j?�S�Ĵ|���j�z�\���X0��C���a[�6��Ư������#1#V���g�r}���)�z��HBzAC�Ȝ��{���up-!`PpW���I���*jhf� �_�L<��xP�߆k��x�+xU�ZU`�o��QBؑ\II��:���L���"L�[X��F����*��m<n�<�(��C�߷lΈ��)���2'���6����{���h��@�GJ� ���6�%�K���C��2�2\%`��ҕe�����6��]mr��?�NR���g{HG294�jX�>�J�r��<b���w��F6�eR@~��y~ <{L��v���yN�p�x&Z��0F�J&�1)VsP�4K�p��pڱ_onY[�߽�*h��S��ߏSuv����?/���*���*�8�GwEm~|z2�]X��!|n�F�4�|�K	rb�!uE~Z*�h̤���_�9����7J�= ��ȥI�Vʱ}��:I�M�I7L���H6����+*���B��88�܂�.��&dh+|����ne�d�{#)y��E	�&�[T�װ�<�w<�����ߏ1d1>�ȥ���>�ְ�g�3?+Q�*� ��67�o)Q����V^��u+b�����<�#E�����������l�F�ѓ�[5�HNraո�4����x
��/�3�suu���Ω�m�
5��C��z;����)�L���u��c0N��1�#Ǜ����Ĵe�N�R(&q����NB�r��&�BIX�;�1�:C7�	桥�����+��K\��p&+���/��'��-s錎��9�"����iF�"bc°���4L�k/�x�D�j'yۅ���1����_�R<�˷�Cj�%�QL�*IS��p̀�Pv�����QO!Nt���tw�/IE"����������H�H����&�g����EM
��XX~�vW��t�5��l<=�ԫ)ޫ Ȃ���b��T����X��U������ #
���T$Au�����xs���9�3A�|�Ҕ%.tޓJ�L�O�V���f�^�c�%�19�?=���$�y�5�����Ï���
�i�c�0I9X��h��Eԭ�O�f�:�6x���2��ܧ�:�ad�'1� ~�^R�_>�<�*�R`χ�
uF�����}L¬�:S�����|y�:Mz�`��ud���0�XO�*74f��;�a��P߱�|]	��_�����(t�t��_��z��W��I�Dg(i��2�����&��+�.��j����G���uP7h�Y��w>[�R��;g�ڰ��gi�heP���m��~��b��6g
�?�+AWW��8���p���S��Ç�3�{T�G�Ʋ;-_��/�Bw%Ƿպ#)�_*=]�kÚl����r#��A��ռ�"`eԛt�2��/u�U�?kh3�T�qmHB�1���c��Fp���f>�q1->����k�W�����tD�V���
	���⒩���&�c��K�ْ��;^��{��A5M��s��mI��e�!�O��ɍX��<-Z�h���4$�@i��NNsI������r/��e]ǒ,�T�[����d_��K �Y��?"�E	�#F fVd*��8+�~g5+�|R�6o[�r5!xG����9W?��@hᆧV���9:l4���b���r��������1�nsx�wA�Z�����Lx��P-:��	��҆,�p�~wP����²U��kE����.���t�,���^3-v9�bP:PO��!q�F�+��PZ}àP��]�^��;E:�������\u]l\"?^�7�k9�i���N5i�U�<r_(�ݗ���M��Wq�W��&��?)Ӊ�} ��7��Ƿ�Ry����H���䔢�����4c��~��<���<,�b���;�L�3~Z17Q�.�M�8hy^r�R!f<�s2��`%�UBRѫI�q��,c��Γ�o��ҟ�e4<��`F�M2Pܽ�9Fzw�� 	p0��?/0�*Qm�P�CD�*�vp�^Jp ūB�<�y�xҔK��h�)��'\}�� 5��L�街w�Y����/3N|.Z���G�gI��y�Tf�MA|�� gt�̬�·.���ټ��0�L����.\��8g��#�4�W �щO���~$�9s_�K�{����c�ɞ��=Ft_x����aUX;�4��al�i��JĐXT�p+��I��b}�$~ứO�X��#}�2xSw���1,���p���:�ԣ0Y����fLבW��ϗy [9��-�	/��4e�=�d㈡�<5��J�3ޅ��.�x��
�-l'�/)pn��t��{n��	Qw�	�a}7�s�z(��hx���I�+H��T���Y�����&\1��b�h�=�	�xɽO(|яS�Q�3}|��\����wk$4���a�1/7��N8���an	�3�Ҟ}��e>�2�T��;3Zy�ꦾyy��7�S�o�B�Zp�r�g�l��#�$5��a(�-�P�z�y��z�,�&��b�f�_���e�h������C&�d�e�RY������
������r|��mg���'��Q �b����.���.hZ��=�F��H�!	��Rɼ&z��N�pȶb�����s����1+|�d�F�ϲ��dU���k�Sm|���M�:�G��5 \����>�xu:#dzC)p8���sN����xmO�{=��a�	h� F�P:��.��7e��G5vO�#D� ~���Y�j�V���m�Ado~�a�7��8#A��������x"G+����i�����*�՗ެcwf;f�z\����AIbuP7���u�!P=�Ѽ�^�.���n����j�ە=�`�W�p���N�,V�8��7��� j�п��y�������k}���*��t{Ͱe�A��O���2O7�=�P��E�*-x�m�z�)� {dh[�����V��$���k�@+������%�~C�X�Zs�� 6���V�=�2W .Y�D=?����rXA�����ns6��4��x�N���\sCmL��%�@��h�i^r�ϑ�����=��)�ra@��@#"?��~7�G)-�q?Ԗߛw�gf3��~���%��TY�xW�uǿd��3� fT��g��/�?��K`̛���쾆X�C>Ld��w�Ha<�!���Y���n��_@i\|�W5�����2�il몂!�dmy6ɌX1�of��O+��\��w$�m��(�8�M[����Kꭊ������*w��,�2=�PY©�bF���\����O cg,��蓸dR1t� �ᮞ��
��N�����'r]�"RK�������=)hx. D�R7l����VS����!6��߹�������?�`R�B�Ň+펅!��ȝ$����\����Q6E�B,d�+U��"�{�T �؂4���j�f�9�G%S���a��Y9�'�ۋ)q��>�\a�9fcx2D-1l������~�'6�*�zr�,|&��Ձ�g�)��CX�w�����	�?�NF�1��Dv�!;��D�0gb��U�Sd�+]{Fc0���jςLG�I�?��[�[J�`[��@<5��q�����k�"B�V���h �� ��\U�e�'�|���t�����|�P��Њ�ES+�J�E;o��6�p��E5c�<�9��!��r&�K0������8ӂQ��ͱ�F���`[�W��\xb�p�Z*}�FQۉ����Y�s� 2������Є�������,9k��]L�����o�+*&|�/��wn��ָ���,��_��_xPP��_0,�!�+�u��й:
ns�ߜa-aF!�k��ID.n�LT��N	?wm���$��-l�I���n�4�G���:G��A<m�K�k���|{<����Gl����GƳ$���Alq����h+\��9�m7���؉�_�o�����o�e�-���]@��Ig����Z.	`O]TB�wOGFsFZxw�Q,I@ A��4�ǝ�b��#�>M�������G{������,�#�U�O;�9ϒ�Sj����+�K0�Yp#�Ax�c����mS[Jn7�ۚ��,�w�0|��eFE=0,8wQM����' ��O���3�jZ�Ǹ|zӗf2WRr�E�|m5���O��Ta���8��C���=2����,xKNDS��N���@�#q�{�����B���,��-�z��3!�Y��(�I�3/BI���vZ�V�3�#^߃;|B��	�Ӂ��q��<��OTjb C���%{?.����\7]z2?�!m��x*ϭe�����;;%����]^�$��+��%g�]t�ʏ�Q�sP
���kw6��«}=�Q����?}	�~'8��.�g`O��[������'4ȧ�V Jcx��զjsiF�U�<�?�Ɓ���ChH�mָ�@y���VR����M�x��+ݗN�����W�y�]��.��'\��̽�C�cnX��JW����-��K#K|%�[�w�{��p��� �I��P�����%���L�[4cF�.�)�cj�P0�Kr��v`謄�����=���t�y��Vw<�kѱ3R9����|��q�|�` ��#�ow�
��W9!�-�%�R�|o�M�U�.�����܂u�̀���Z��djK���9(��"���) K{��9�3����r8;����kn���Ƌ�L�;�g7�w�i\�;vyŅ��mv�~0UY~��(~k�W�8�؍�F�7��[`�T6쯍!�-�`�(���>&	D��eK�<ڭ�;�_�������_�:���]K���zz��m��Kzڲ���g@t	��,��wN �Q���Z�1Zmń��"��HB��d�>���q�	?h�L�����0! �8�Hꂖ3�����T!�	�=�=�s+�21	P�i�4#�¦�sڛ]�r�m��T��L�U�D��*V�r<{y���o"��f�a���L���c ���ʌ�j�����,�#�?�FU��X{�<��z��Ǝ��L�~I}��~�7�b���&�I�'���n'f�[]2
ܷ��k�w�V�+ry��΍`��٭�	ɸ0$y4o�8��(�}�z�#�v������̟���q;�ɉ�s�&�z�����4�k�P0�j�>O���c�s���[lЩ|�aH�_��a���k8:�%W�Q��^�I?�{
K���!@�e)d�U2�l�W������YRi�XB��ɰN8�����$׮�~r*r-I뫲R*�/�d��)˞��W�)q�י�Aɽ�]L�'{o3���S`�I�Ӈ����$f��ߴ�[b&W�XW&C�yúw�P?>�N��If����9�$�=�n}��%$C�V��A2���Y��2@����8v�B��6�0:�.�bhK��=�?��~���$�1%-:YW���a+�љH;`��Ok{��hbl�1x	p��+�� O��"4J�Y�_��Y�Ǌ�t��*�Y����s}r�]3�_ׄ�E�r���{X�;IC�Y�_|I%� �=�<p�X[/T�B����H�<+ąS�D��,��9���PjS& hB�0>�cu8E�����J�ZIԼlc�8_m����W*j������z&�� �I#Չ@�d���6�=��\N���S~�7:�)�i�L]����<�z��3�%�e�Zk���g$�RY}�ۊO4#]�8�����;N����2�K��>���覿�9E��T�xhjػ?��	{�Y��u�:*��O�*U�̈�<�)V��!7~��|:�m�KM6���}ZfF)R?�3x�"��(�Z͢�(�d�Lᦙ��r].����j�P��e�C�r����k��\47B����E�ѱ՛�$�^����J�iDf��ֿ�������T�pj'�q�^��"�F�gb���AA�أ�#��GLTlF�n�L�϶(����hY�p��t�i��:<^'�|#Z�[3����3�f��-�]��c�bcv��Վ�{c�w�D\�ftoX�M�@��S���.ꨒ�
�'0�v ��j$��X.�m���ʇ7$�x���^R��k�
tN:&!����D|ڊ�i7��H��<T�\��S�imi���8�_�N�j��}�@m~��V�A�Oea��Zu�O��$APe>�����Fm���hU�+�������י���̻/���s	����|֍Z��lD~���*1���|kGBS��8�8�q�`7>Un/'
V޿Qo�_f~h���o��o�Ǔ��,�$�|��Y�pO�ّ�=e���ײ��Wc� @;��|��s=���po�Sh�ն�=N��a��>~��C#�J�{����V@c�FE�(A�j�R��<N�|5O9���c����������wĮF"�������)������يO�6���1�}� ).��F��u��+���j8�Y�=��-r$�ܢ���
�����|k�.XSZ�� ���M��4��!���R�%��"w,�� 7Z�S��2��w�K=C~a��N����9�p�/�;Z�����|HX��X��&��h��vQM���'1��/�|F��K.�6��������t�������_t_�'#:���m�pN~�㧑��������J��0Y�!v?L��x��"��&����!�k���f�a�\;I�	��t�g��*rź��}맦�k��vJ��(����s�ee޼^y���2���f
3�"���Բ�w8U������\_9E�$E/���3V���� ����f��'X�lۂ��0�,�cZ���E��'���[�b4��u�6g���c�@ �'�Q����i|��`}BZ��}2| ?+|�����K�R^�0a<�҇�<��w!�԰�?�J�t����>ٸ|k^��^�8�Ur��"�9<��f6��g��f ��
A��H�m'���G�AM����mg��~&���M���)����&�|]��ez�]Z1�)���������iUC�IPS�)|����'�F�>J���êq1.���Dn����,o�^?������W��K�읍]��>Z�&�8TQi�$&X'��3�7�ak�AS����u&)�ZE��NW�)b��a�Y�J�r��zy��K������w���|���Bk���5�!k��O�#��/6A��!���H�~��qo<���,wX���S��V����K�#�ە4T�a��)_O��9GsM?�����e��`!��<ާ���M�A��u��^'��i�d�U�x��u����ᣟ�����tQ`�Ż~_����.�_Oy�����i�������_Jy��?u]��ν�Z��;݂V��Ȅ�k$֨m?����PaN.���(��q؁�����M4K�4��e���d���A-*���a��P,�)���	�H�Cd)��J�g�mY �]�pD��1b/c�,�b��.�Q�=����N��4�% �l�>{�
�d���F�'TC�d���((%E{ڜ푏�(ҳ��>^�a�E��� �}d��j����"����ŪuFs�uX�B�A����PiUO���Z�Y�w��O~��$q�QI��A� �܊��r�� ��	}��U��	�CSo+ 8E0@n�-#X[1T��S��EQGfLPY�R���x^N7$\�҅�i'Bt[&�H�F�hg�V3�U�+}����UP���n5�76%t�Z]�@Y�EP����Oז���)&ّzA$:�r��I�W�x�(KRS�lh�~Q�I-�B���D5=Z�����S��l�'
ʆǠ�}���������O_�~{'r���o�� w�f�bRi���AH�"���ޘ�-��:m��f�% 1B�x*V��U���tm{z]Ē���t˒c���J.Nw��_�� �ʭ��7���7��@�[�|ʾsv#0<��:�G	�)z�;�~��Z�fl�؏���������Ĉ�u��U�0w�#������T�����G�4.�n���(���i���V�OÀ��aIRj'���kv��	Qt�?)�
U�gReHF�t�hW�&��rG�KBq*��̮-��]�&��e�Rh�X��>��5�Y�֚�K[s�?��u{D��(@�/r�w^H�E��;0"?.�^Jޕ-�U�Q&u��'։:�*�U����ū��u�x6-X,ěG�"�d�M9i�撒��h-���iqiW�WmVs���~��5'�e�}��/���Z�O��Qpps�*cZs�s2x����F�����������Z�U&����������#)b"��>�G��R�SN 0�]7�����WJ���2�����.���/[�'f!+ֿ�HJ�N�!�cn���]�e��v��zN�i����dNq(+r���Z��ũ'!7�M�槹M�1�h�c���Sl�ki:bJ j|F���z�m���IJw��`*��Wc��F�2%wFlյ�:�b�~��K6J��̸F7]=�FMm�,mn��'QP2&�����4��AB�����b���/�q�xU0��6��hx�n3H-�c�=�4��%mc9�w��rF^���O	����z&o,�&z���P�K�}����c�^R�7Ai��y4م���y4.tm~�Ý�ڪ6{�6�^&"�G��ͷc�%^K�Eǰ�ح���mO����V>�A�B�ZY��5\��4])��.l���Y�
J��8Ҳ�^+�#�xV��4E�x�Ý8�ab=Me���Kǒ5�bi�;�,���뉔L]ʾ�H�?Pk+��G����Ň2����xɃt8��#�:�Σ�ZiԼ��7F��(�-Z='�V�"�r�����P�Wc������tC`��c�9�і4xG',j���d�5Nl�����ZLƏSG�AiD:�*�&]f�Y����#����������E�#�}��"��f�G�Vm�,�i
E�aaI����%Uq_������#h�ӄǃ�Юz`��4F�k�[��I��6�er�P�V^\_�ν(!kU�Pt�w��cD�������3`��{TD�C-���scU�^��o3f�+��ߥ�E�^	l� �cס���G�v#����Q�	羅fG��MVw���ýT& ��}�{�h$)^����_�@f��l��l���$�:.�G�÷L*1�lP��DI�%��̨��)Ï��훎D�b�).��`W���1s1s�'�"+���k���{��W�w���ꍢ�����k��P;oTn�g�����R�������|౛�f;��k~����k*�Eo��8(�B-?�?��p���zhA�Ͽ�s/]��h�˺c���D$<��}��غr9_Cne��a�'���D��c�_��ST3�C��h���k����}�#K��c�w!y_����~I�)��k[����Z%��.������<�����0GΈ�=2����@ܞ�S��U,�����!6�o"��]���!�%�?3�s���p�I�wz"B� z@jD��Q�o7Ok��9,-��Ԗ�d��;I�ǆB�9����wc	 %�޹\S��]���]})MLW5��LOĞb���jSV��h$��)/�~.����x��*_6,E�{"ɺ/��2cvQAt<����:��#��xp뒙��ZK�p���럎$��O1��Y/�
�B	/����<���=�h���xܞ���EZ���_�n�!��n��S���6<�kR;S/��&�Q��z֥�����}�r/C>K6����+�����,4�����X��U���x�mN�`ѳtrwG^�rٚ*����QN#�ͺ�#����H��}��&~�d�Д�OJ-,h�p�HX��z�AH��� �}�}�oOU*E@���	�Q�ᯁ=v�'�)��zwiuu-��q�e��+"� ���EEС1m�nB{�nT��*
3xɎ�j�[z�	�Gؓ,���=F \�K�i��$�]:0��u�Y���*x���6�D�B�ΐ���
�@�fs8}7&]H��]?|� UW���ۦ�������iO�<|>��¹�� s�R��)�Yì�.0�[KU������Fe�9wIgo3�|��,�)w�1�y��������TL���Rq,��F�a��A<��Q��9ʙx۱}�Â�-J��(�9]�5�wgp!���(��d�k�(k
i�';��"�����[�v�q���dO�[k{��& �&"���\�`{}�pa��`-���[� ��nt�}� ?������wi(��Z�v�I�x��P��I��uLGK�+�l�/����$�=����j�mZM�Hj[�����);��2���m�l�"���L�g)S�3���h
F��Z,FѺ�/L���X����}�~�<#�9��B�J���Y飖\w��x�:�َ'���;�bO�|��K���E��؉Ť����
(J"���h�)�<���yog�%�ش�:"us?� bD�٢1EB�u^�c7jYjD�O$�{G ���4cJ0^��`'��I5R�zy�w]�d���T�-�]4����,�xK7�P�ޏק�P�z�N�#;v�ʐY'm!�!�^pwҩ3]��"26�����P���eW�B�ŭ7�����.ɹ��%�[Mg����|�g�-��I��_�Q�dg�;�}eY�!���D��YF�|�b쬠�a�U�:��n��͹Nൊ�pT���}.M�\��� 4�ե:�xn������Y�w�\��V�ǿ���`������r��_Fe��tB<> 胅$<h��,$��z�Q�p�7�ψ�F��0�t�.i�S��U��������#��9K,�`.���d���Y�'	|���S�L!��{S-מ��f�
��88!�[Ȇ��3�����bs�Q ,G����_=�[�m����4�4�TRf�}iA�������*���k䢍�5#�m0�Z��SS{;�-�~�2��G�Ujiv*�}#6���_�m��>9m�
�iߐ^��@ � g�V%�G���k�q�	 [a�B-���<&m����n��>�l,����n	�o����.+�ӗ{�KN� c�x:����u �c�\�`��U�m�2�H��ܬ�]O)��G��K2i�!m�-�݊F�T���6IO%<;ҷr7��^��O�}��>���tfÇ��'j�i>��������Bq^�`Ś^���Hd�?��mO�P���X�Tg�+$r�'�n[F]�z�*�I�z�
>��CSVG�nMD�CW���.��1�i�w���r�s�ɖ<��DR���
#�Ǵ��z��X���b���e��xd�|�_��z�l�ÆZuC,�K���S�a씇_7�,�Y�/}��p�;���r�o�g�sNҩ��ѩ�5�@����T>�.y�xY7K��1�N�b�#�\-~��z?Yg����Ғ�7�?��76_#{�t��QH�;�4���d��?�;�%n�n�G��S�ʽ����`'��x�C�	S�Ė�~Jn��!@>�#=��}$&�Z�#<eY�5���|�q�&�^t�F^S4H4(`��KY����W�S��qn��`�320)	~��]�1��o�x�ǹ��U�L���/�@ˁ��J�=`&E��q���9�붩d�xD	�-�?T���Z���&�G��RO`��м�{�`��Vˑ������N	�]F�*�܃���rj��n�A^�ϋ7=�N����RP��I˃��������Z[}��XJ8Z�H�	�� _.Y:�)^�(ㆂ���S�:WO��F���|�Ϋ�;������⸼Ƴ�I�$��O�"�Nk������MB�̄����l�[:�A������eCd.B�c��SO�8J�`UPBCYl8[%[( b��[Ú��ݶ��ծ����}��Hч���a�ʷ����Q���|�^�\�C������+!%Xx~��������awF�#�w���?����`�/��i�������H]��J���e���h�#_C��j(
��氾�F��a�_����APn�7!nsE�E��[1[�Ĭ���w$��j#�>�c<�Zc&�9���W����,�3�p�s�<AIsΔo�ӎ?W��Su<�p�Ac��M;��~ ��Je{�!������m�qI�[�k>���V����g��)NK�9���8q�$���:	m>+1����p5�j]$�!�c-0��x�e_�񘴐�^hS�H��뻧	ZB�#W܂�FiȆ�����X�'��`X���6-D]2wӏ��ϱ�Q��=�f������}�u������& 	��7��͜ثMg<&w���>�EvD�����ꋁ���2E>��Z������[���T�K���X�fX2O�5>4�dx?䨷G���a���&��A��"����J|����5�,#����a�|�T��[��P�y�����Z���c;u������5����U�zW�/<�[�+�V���*_w��1���jԳ�k��|{��Y�U�D����`�������f�����(��c���Je@��=�=��]<���;R��WAf��l��X^	�9#����1>�Ԇ�o�~�&tf]��N�U��ُ�׽�$��\4׋��YM�̩� "o�<�bI��^��Ɯ\�\Ө��m�-�׵��s�*CL���4��f�5�E�i�8�E��_�{��&��`�����>`��A���A��H�9��^��N���B�Z|-�ia�\��30Ks_/�v|��s��)�@`�0]�۪6�o�����n�D������0�,���s��+9�1�;�U줥[w���V�ZΥ�Ftem��+�y0�7�?����E��&(��cހ��Q�d*��o>��v��
�8j}uK��ލʗ'��#P*Ǖ�c~wB��:�MߚQ!f��������u�>�&~�u51���� ����z��dYM*��0��P���_X�����3.����e��>Y��c�秳��5& �uZ���5���F��o���Z��E�V@]!�C8��4;���`Y���ѣ��uЩG���:q�Z���#$ԏ�U��J��tvc�&���I���H��7�Caf�j<�#e\sVv$t��	�^^H�PWbe>}���Lé����@�*iN6�Ә,&Z:~��Ć��E�T��f���	�� �7��Wt�E<���@L�>-@{����9�F6��>3�4v8�IP:.����<G"������*�?ߟ�����`ilk	�����I^zV'�:{���0�U3�}�4Po���k�BlP�+���gjF���M��땜W�z��ɦ��ܙ!j�Tt�^�5�45��tֶ��I��/��:�* ��T{3���R�@X�[�Q��I2nIp�Bc�[׶g�gy��lhB����3�wQ����(��R�'8��x�7�?_�(fD$�����-+��������Q 0�\��!�]$}�ۗ(k[֊?��&���(rz��y�z�r���dN�5�d�zj�<�|м&ك.��"�.��ȕhX���g��ԁ��T?UrxdCYX��D��U�M�t�̚�����Ï'��&Qӌ���x�v7R1�"n>1RW{�K3�{����S��M
�Q����eӃ���y��fO�J�9��I` t��&B�Z���*c�U�Y������Y�ٲ*\E���d�����<�\u�I(^f�{��o��t�\l�?��e�x'�ayΔq�h�����M�,ޚ8�;��'�'EP� ͵�I���1����(��Q�塁?�؏�Dȴ�9#��}�u�_+�R�қ�e~3 $�ɺ�&5?l
Aй4=E_n�k���Pܓo�I�,��z�{VM��#���:t�����3���'	���f���Ƌ��0�'ƫO�ͥq��p�fY��8}�����{���yT��zP�[OK�{**� �Z��
ʙUڹ^+�F�I��z3[:8�[EYz��Lo�M�s�&�[ĉ�FL.�	�)���Ѭu\#���.]-^�*5~ z��d����\���vx�r�m���eJD(x[��f�sl�V�(�"��m%��S��tm��o�	U�0	7�曬a�EI/cŧ�>< ��f�%"|�e��[�w�����GA�\�9z�;��#�Jr�3ż0�h�����ѫ�m�
�e�%�W1	�V��6�c��*c�]��k�i��9ѣ��X����%�Ӆ[�+' �7<^S�Np�%R�����2�58o��W3�<X�e�1E}��Mg����X���w��>9]&��җ����v�=�Qn�b��4	1��+��� ����k�oQ�� e�
��-�T\n��d@�AO���5"S����W��!��3\s%Y�\�o�pm}0x���^l9Mn��Jj5�0q������
]�Rl��=Z��M�h'�U>��?wyg�lp �f�"�C�p0|���@w�'���W�ĢU����H M�������"�c������E^�ׇɤ��֖��ˎ�Ǖ�9P#�#l�d%'+a/�h#iE~�P�bc�h?n�8����\���x��O�Y岍��`W�!$X�5�"|OMRt3d.g��:�~�d/���LG����2t�8]�aβ�Q(��a[�x�����/d��aZ ��Ω���J��gm�B�j������6�����@]3�Ka�P��A1���T\�]Jߝ�l �p'(O��n�҉w��+�!��k�FF��Z��br��j�)��P��'9����.mv��6;�����غv�t.��Z��.97�hi��[���XҦR?8��qdt�x{�0A����w6]i�J�Thr����PIh����%�(�5ڂX�-�$��z�@��z��ζ��Z�L}k;�Hv�:}~#����tڔ�^��3�\ߠ����~���H���C�����Y���=*����ݰ'g��/���gUJep��;����X�qG�3�[��O��ꤶ�[���L3t�I;��'*0Fߑ�lO�-i8e�?1��=q�M�#��q�����Jo����ΪPO��$��|mV2G,����8���GI��P6��N�]: !]	�}�Zw����ibZ&��O�T���H�vI���J��[o����[�|	(<����¦>��-�C�G<ӯ�T�VS��0U^{�CA�W����/�l�KZ���4�\�E��	>\I��f�	Z����6�߭��ר����A�c�Mz$Q�,�=�p�n/�iRȭ7-1�TW��,c�ݳ3��O^�����c��ݚ�zZ���{���J#�7�"i�f'<���H�KVӆ~ ͍>�tǅ:��)��f7���������G����쑘��#��(ԎE�u�^0Ň>��Ф-D���d�W��~�ն0)�t�Y��mړM�Zl�P�]y��]���N=M���y��?VA�9de��w����ʀe�|&Ϯ�΅�/���Ss�M���Tj����qښ�-��%l���D>����e��`���x��J�
G�ӹ���7<F�6_	a��JH�e͉�F�����dt�~����U���|�h��g��[�a�dyq@=��,y3���J�(�|T�B�����G��VO��f(�劑�9�TA�{U�hf��{����D���`w�e���)m�s>�@}�P��g��1��D�pn&��%.�n����P�b� �h�(ǉf��(��}}�a|9ѻʓCܑ�-iqd�[L�쯄�\gPJ�#�&;�m��V3��ގ�"Xۿ���ĖtV��i|(�.�v!��Q^o?�ԕ�5V] z�þr��;��I�V��R
&3"�Djh�P`䭱���} q�$sU�=.�.��k�1��^%�w���>�� �V�~
Vs��?����<X�u�=�ܼn�%���f.����I���	VBxi�I�<�i��"�F45��3��`r�vD��Ub*c8e7-9�Ał�A�2���#�pgij	�3ǜX#��0��&���)��e����S`�MԺz����n���I�@�
ᄌ�L�5T�[����uO�ޟ��[�iͥ +(��㿵��y��/I�L��=y\��vIr�^(-�p����Zu,	L��s戍�;���\II)ʭR����xj7Ik�i�/��ϑ�$&�WO���>6�yB�eڒ1j��5���_��6x{N��{U��f-����%������e�D�w�|��'�a���j���K��L�O��ĩy��;9I]�@�.�H%��9\�����]y~�\�p"e��=1��K�c�.�j1G8��&"���e6�I��8)e3W����ۄ8Bм�v��Hb|�u0ǵ:|��)���f���	B.���Ŷ�Ĭ�n�Uti��l�G�^�
�+���h���
v����"l֎��f0s<*�Ѫ�S� *�����)P�QQ��a�I.a�p~K�tS���+:r�������ǣLӫ�Vß��_
-;U�yoH�s5=�[��ȥ���50�I-tᗭ��2;�;ʆ�1��W�A�[Y���O)J�S��FT�gb6}�r�@�:�t	4ӆ�ۉ�v�Z�Y����$�7��H��,���7��<�°"���\�:B�,`���s�K#q.�� v�zq�q�S�#8j���3�x���W�AmZ�N��N�1n���"���P#ē��֍���\�}�x�,u���mV���K�����a|�~�㛭�]�n1�%6.a����M_��%�3��b���t�xm\��h���%*�!A�x9j��z����"��XW�A���#'��~}���|� Co��8�9�E���m�������~'�ˮ�-��E���o[�O8;
!�:E�@��`ڱ�]�3tw�w0R�p�c2��k������m�|�U�J����0.��wQ��6;���zs��0[�ŧA<����Y�Uò�d;��8����-�����gc�������x��Jm%��-�|����cVsq��4�}�׭/[�o��o���r���j����iq��;�׼��u���vd�M��[��1m�Tk���,d�K{�>ѭ(�z�����Q�0jl�`"J����Y���N���Hډ����@�2ZĒ�	=�lhf�ըQ�xSX���͸K�IוZ�,��1����i�W��8��4��{	Ū=j�ic�4��K=�7���1>�{$�2��̘P�\�������*����WU.l�Ad�_���y�X���b5���+5�+
���g�_W�H�����TF���%��2��P�!떢� ��}�C�Ww�~:zS^�A�j��-���Z�V�zo�j�"|�E���"�g��4>��_'��B���}f~�5dKv+YDҁ��m��/�\�c~5'���ݰ6��oCإGlz���Z��H��� J�̀�"n8�ԖL���L<�����d���z2����!%�F�P�i�(�,�r-�ƮHyO�_Ӛ
��C���
�æ�J���:@�q��(�z��!��>M���:a��
8Y>FX�.��P1��Xϣҗ�m�u��xG�́�{�(�pfy�A~��������}�ҟn>z�}��x6>�1��`Zֳ�����GK�z�c�4��Bj�k;����QK��
��e�!pY�����Ud�����1T�4"W{C��E;�=������X�=������h�4u9�C^�a�À�`.`LbQ���:O`��5��ۻC	$.3�.����y�C�Q(�U�r�}aU�6���5�Ï-�`�"��F73�8����-��q?^�xl���Pv�֤)z½t`j���X���gm�1��q�zv?/�T�Z��3���u��qi��a5�`�Hc(�9@�����*֖�`���V�����Y�)%�zYkcZ�[��w���+¥���.���[b��,��}}�2�]�Z*�\�h�V��MK�_�����TE/A5�����D/}��ޣAƁLy�6{3D�R.�����雰O���v�Ýӆ�'$�\��'h���a����q���WA N/��m�����D*�}�A�O�<�C::6M؟[u}�f�:�3W�_%����>~���*f�����WҖ�L��a�_�wk/��_���;��9�)�,��jKP���P����Z�l��؊Tu��轧^EM4�a|�
�"����-���s�c�)YR��頝+{���w�$��3����L5�0=��4�O��w�gǦ�i�(JX���3D�5�[�"k�q��.y�!InB����.�������D(A�����
xQL���W1D ������w�q'���$�>�B�����Ĵ�3`��c�Z��9ĵ���������*T��R�!�zr�/���� �'�5��v�0���]V�7��H'���:۫�韰���E�Ls�/��F�qW��@L��!�,�2d�6[Qr��7cr&�vu�!�@s��zU$͐';4q��]�����};N������xtVJ�M��k��H�[������HM�(D��,O�@R�X�~�nJY��yM4���2J����2�M��ŭfWY��!�^H�
��`�9{Ў�����h{n\<�P�����/�o 0�8ĕ�B���I�i�1��|�?�&�/咠�x�-vTzr���^ ��\ʁ�����rA:�r�I�|��tχ/;��$j��V<5ᐘ����=�F�:<�2ҁ0��U%�0�m��p�X�갨@�cver�d��F�]c��04��LR���Z.�������]��Y7j+7V�|ֆo�N;������;�qyNC�(_�u�� ��@N[�_7����%m����u��Ĵ�$��.�,=��3f�P����+�uy��5��q��l&:�U$����9�ed�80y����5��~��J�فO����(>�!l�>�{�Ƃ��`������������ǉ�׶�V�7��CAG���.:]��jAt�Ɵ�]z�bD�=;�f�Y�}�� ��`�ڸ�o���;�R��ԧ�@C��l���ߕ���0�|�g��Z-E�U��Ԇ�@�s�L��Kc��('�1���3x�7'`"'�xdr�L��-���g�1� �uc��|�9E"�y[M"=�9yC�O������5H�y[ФAH]]�{ ��02�BݫW��<OABod5�Q�?�w�����[�c���؜7�V�	F��b�ّ:B��A���\u�Mfkd��@/3���~��.�C��]y:Y�`Ѭd�+~����	�bR�եR��g�e� M���� ���p'�6�DL�RP�[F{>"1�ʪ���@��;������ʢ�F�v"�v�Ta�����p����숈���󶚟�y����s��-@����X�� �{!�Љ�Z^��z���wJ�X� �A�8��ji�}������Dz,���22��yy���ڇ�r��[�f���%7+�Ĝ5��A��&���D?��Cj�x�H���9�OG�%"�@�,Y������1�`.�7������H��-�q2!���k�Q�\C~.0��YϨ���϶N�6����^Ժԃ$��;��]4� ����ēba&[���n?@
*7`�!�ݶ�
b"�H��e]�
c�6Ia��ʗ�B����^!�	�9f����5����0C��"Y��]ߑ�F3�p���ڼ��#�^ntl�{fB��Y�EU/�ݕ��R[�Q֙�(I�����`c����m�H��h�:jo�s��B�'�؇!><����E1�F>���N���-.�	��۔�%���/&��Ͽ�˔��dօ?�I���܀�F���_�L���t��>HG$��H��?f�\��f޸��?��ҥ���Fߎ�h*�zT�����م��0��:?�eٶ�����CN��}�l�E����w�_StJ*|Yu$����ǈ�[n�?��`X���b�V'��጑�uTm�L?/
Բ \>4.j#"���i�^A�f���ɘY{��j<�jű�'S�P}��:�3����W�2�0�)o�zeG"�ZO�'^�ʺ�y(�z��A�����^��oA�I��������=E� �>��p�fV�Vbm�A�'>Ӆ3�2g��Y\�Ԡn1<��w�&�g�$�?BXP�	Hݶ��kvꔐ�#��+�ָT9e�~��R[�I�T�V��Kx��:�N��J�����M�w�N��{�v��+l��̻��^ˬWR?�b�<�P~EŰ��Y�:���5J�N��9T"h����I�y���U���3p�#r`��>
�#g$���Rh�H��	�������E6+1�ص�1�����<�)=�V-��=~8�OC��80��YE�讨�c�J��o8I|�Ȫ��s]�c��)JL�#�U� ����J@|�Y���ϵ�S
@c��ۑ.IjW�7@}�QÎ�q���d���F5���o�9�sDAs���YfC�M�^bNf�4U��N�:9ѥ��������V�ӈn��x^\a� �n>�n��B�3�x1�2�d��/4�F���.#µ;�j��˔�}0��K��!��|�ڭ�7�ձ��J��C0d���;�$UޕQ:����"�Z-�|���|nD�,.��[B�A�ݔ2k��*/ʻ�k�2��3�lM��ҫ#$Gt� ��g�L!��E�|lp�F�;�VA��yt�ic� gS�p�-��y�8x?�S��o1�Ýӵ���&�`fC
s����GEsW�����(�g���=Ŷ�I�P2)��y��B���"�@�wJ_N��^�*صr���}%b�M���$�clԂ�@\(Լ�@C����Gڬ)Ƃ&ҟ<b*��
�
i�87ܔ~_�c+lJ[���K�.�Ẇ�8'Ǡ�~���[8�)���&Q�s8ԩ�ih����Zb5)�b��^͸���F^ �"��?��8���y�a��Y�O����;R��&}�P;��F[ �<�"��*��m���7X���Q��z%Eˊ��$ 4+3���9y\����ó�,�
+Q�=���x�����-��$�x���!�1�ټ%"�6��"�����3aS~��3je;�L�-���ߣ���8���0�\Ǻ�lv�u���$L�[��jc�=R��Q�+5V� _g���+��A�S�t��l8t7I!�`
o
?j�HiM�|�=@��W��&����
%��n��[Ѫ�L�ҝ2�e0Rc���L�\�^��LM!0g��|J��ʍ�):|�(�K�<���T�g�%���ʞ%�������bt'���C��q#��tF�E���<�+.��(5�H`�@�h��oǿ1[�j������,�!􊝗��[D#$�p�Ol�C�+^AT3e��qg��Et��}w'��,��|���y�@/>�S7���[�d���)���-�_v�W��[�J�q���(�%5h%t�D$�Ho�t��hU��Z@�L���^�/��+4,~�+%=�ǧ_\)�ȍ�K;��[�
�3����Xx�(Q#+n'��w�CHA�����τ(x��k'�P��Գw��L8p�7����Ϊ�}��%U�����{x����L
�j5�A�OT�a�y3C����pj'i(�ߑݾ�	$q0z)����~�=�[i^����M���a�hz���`���g����,@���	� ���%��a��"#Ϳ�Օz\5�VP
�q�W$�:�����`��K�ZM8�vi�g�%�!f�-}��O�x� Ε�Ca켢 �� c��4
�ʔY�ޑa0˝��*���>I.k�e�^"���5M��%%s�a����4Y��)θdb�W[V�����-kA�v���ODJ�q+��BO��ku��&-?�;#�2{��po�Ju��V��'�࡭G<�}���w*;����xG$��3���hq���c����V�0h�����b�>�룵HøY�������'�i�]׽�'�\Wd��ò�A����g�R�B�H��y8�E!y�G����|�j��:�H8���RA3C�t%��F_�7�Y,)��t�28P҉ll~��[�َ��p�.��v�k |a��*��\��������l��>A��$�38�ҝ/��$��Ѥ�'�C������
C�x��:[ 7�v����V�F8O&Q��v���"ܟ�0�ԥB����b�-��k��0��f,�?�հ�̐&��t%@Dܱ�\�]�
�yw�9�?0�<|�ʖp�ups}���I���E��C����T�Tp�Ox�H�5^3=�%�e-�PA�q3C�|ؗ�������S�\�Zu�?�w}��Ym�tG�d���-{&$/��ɾE�TO���؛����,+���y:xt<���m� �0��D���D;�S����aZ�O>��Z����p��B`��f;��M�(<ɵZ��4Z &0Q�k[��q�k������
v!�L)��1k4�R^�n�ˎc��z4��0l�?1��F���`X{ۅ\Z��-�́Ե�KE��/� �!%�����5�%����K�U�J4r��eN�-�ׁ����l�G���rN����K|i'�о����S��A{��)	��>�oCߤ��f��"��V8��c��*������Y�M���^��Ա�bC�[��RVF�1�����>��J��f㽇�|��&Gqx*�+6]����=�1�w�d̠�POv���u;LOd&�)��A��ۿ�L����k�Zk1��?7ż�>��B�:T��&G��w�V�
�q���4uː���c4"��^B�W@�-H��(>�g���:��WlzB�4�Z�au(�\�r���F?�����/َL{��`��]8������=g^��g�^�\�~�����Z,�ൄ\���Ƒ�9CZ^�R`Y�#�[+�O�iey�q��l;3���iG(��ʺso%뷥�Bea�nP�7ƶ�Э	mX�ōOڡ��r9k�}��C����?�W#%���5'm:e��������_�R�� {R�Co��T��3�v��G��y�l`/�1I+G�c���$�����]k<wa?Ȕ�c��I��]�i��X��7�!�WT� {��2Ѣ���ʴ���Њ�Ī,�������M}k��o�1GӬ�p��vQ(Vf�yVy
���pw@ɵ&�\�nOn �Mn/r^��0�x�6�ܶ����ptl�A:��g^����&�@4(�	�Fv�(g�Ӯ(�
�x��jJO2-Mya����[^f��f��b&
��{�u��.�ԏ�)�ۜ�d��Zn��N��Pq����U@mMe$�j2�k�X�/�.��Pn|���`듞�EuPg�ޛq;�έ'"�)n����TgI��Q_�6T�s�pG����L�=|�?MG��
T��+d���]{[\&����r;5�?�"�(��՟u{<>B�w�9��S[�`<���p*�u��Dy�a�y<��enNMň��e��&yf�]A5��[
�ӟ�����V�#�o������$�w��v��_�6=����>� � ɫ.�B_�/��F�(��)�W� ���mD��u�q=/���j����y/g�# 	^8+ip겢���ǂ޷y�*B��o����.�� 7,���C2 Ez7վ/s���I��v�р���ɴr=ȱ��M8W���M���N^���ϟۢ\z�X)�������[��I�qO��P��Jruc$��-�^�1|g���{�c��oƝ�nO��6&�R��F_��u���S�a���u�HW���-Xt>jOn}�0;��fׁ;����7�Iv������gt��� grݎ/(ޯ�վ�E�Y(�9V�A$���V�����_�B�n�Y��P/1���*T�0�Br{���h��r����� ����ݰLj�	��0m`��v�K�����[*�*�l�(;ܼt��ed����o~�^��|�e������&�4+\����QFu=ʩ���X�Qxd�z[�N�T��`��r������JX�µ7��/����FPc�"Xș{0HBm?�n�s(��nyh���U�`I�[�kV5b�O�MHb��w��C�w
q$V���ń�LA<�%�]heq�i���`_[��-զ��d5����@Қ�CLی�B`jkc�¨����<��yxS���rȤ �|V��t�f��j�Byd�m��&h"����D):J���H1\��������N��������mL�l:rP��/�p�D���PCI��F��d`������-�r����	ý�*���Z���
�}�1mc���k�j P�:9����  �7��AS���u���A?'�p4����x�up|-Y<0�^�{�-'dQ$�[r>�.F[`��=UB_��^�q��\%���d����h�n{�o������{->v:�)�ϕ�(���S���S���c��j��w��8����Լ9&$���B
���/���`�C2]8-{tʶPݶ��;zY�Rn]D�%�G��H�m��
Kl(K&�)���L̈́�5L5�B^}/��ӿ�:���	��y����r�2�q�:���k�T��+�	Эք�À�\v�<A�����:�Y����|
�)_sFdǈboYc�e�Z,{$��V�HQ�P��W�$>���)�٪"r9�.���ï��YGn���~���7��*����i�>v���eⵅ%��@�|�e�c��`�aWB�?j��cm�?�d��[֏�f�5�Qlm�/�� 9��?�v��W���t���9:�N9�k����'�� ].����e2B�3ܻ������R9�}�����R} 5�I���L�;0@U�\����h5�}9�x&�8Q�tcw���=}���D� �Q7���ȼ*w�k�G�"�L�Ӻ���^�ߜ���6�)�j %v��M���� ����?H�;�&p�l�Z���zo��F��37f�&� �`y)����;�XR�E�I'�I�Q��P�<Û^v
E|��A�Q3����#:���'D���Zz� qBh�E�����CG����y��9��j\$�꯳ai0���m���`��ݬX��c*���F]�v�¿�U+�MՍ(�H#�3G���簒�����/�O�r6�U%������۞Z�l�h����_k	�o�rZ�X� ��G��^��)2/BN�[WyB[��i/
��E�v�˘��SY9F`X��\&zվ���$^��@��^P<ǿ~�1j�
����A�����3jFL�J��K����0���O���Q�����/��b�`J��D|/�S�PW���9��Ɇ"q�@��6@=�!���v�ߘ�ӳ��ЁY!%I�:�b�G��:>���}-}P��`���O@Q]�9�X����`6�}C�g7�@Y��
>d5�Z��O/&�٭�t��4��j�WS���ڵ��r����U��g�-�[\�����ס�3R��t	JvIO�47k�_K��7t�yg��&�#����N�K�fVLK����\[�����D�
��A3�6�Eo}8A���cU2zF�E�T�C}ԲM=�ȳ�O83 ��4� �P��Tc��Cy~:��z���qF�	�iZ=�J�s�L{�W���W���W|���3k�3�A �-9��e� C���!����ic�O+;t�(8�8�^B]�[HЪ�3ZEv�Iܗ,=�q$������Clh��S���#<cmFS�Tk�#.�e����k�SןՕ�뢂s*����Hs���zG���������"�RVopi2�'XI�/����(�Mp}�H2%1�j�DKؒK[��������y=B�~�o>h��kQ"��[Q%s�/m�M���g�c�/3�/�����R{�+'ʚ|T�SίfR�2�7��"ͩ�ϋ��%�m�>b�a��	�6��J�+Fw{��(K�%S�תfĀ�BE���'1*;��	M��U�s��^hz��1��`�])���\��J�`� W=Uh���>J�ϴ�@ڔ�)C�6D�;���ӷS���%�#�K��[��N#`0��R����A��t-A�@5@7C߰����;�4BbԞ�V��$��:h1�g������V��X�Ά�BR_Φ�$&ڰж�ڹ�s����*R�Oy��P��m��v��-k��3H=�*��<��)�;lv|�Q�0��g��y��K�4'���"`)�y"j'�ʏ��Z?������������iO��#��'�=������C�
�t{���K������l]c$�T�`��������K|*!�TYLzɦiO��)ݣb%�_@ӢW��KF�$Vz�:��S�.�9>J2�(M��'C���`4g]Ɂ�
���
G�/$�F��#���S���Y���W�d�>/F���\=d��z@8��K�L�i-�>�M�)!6�5�w�w����#j�|��3s]gc��qٙ�\�q���,Sm%R�E��'�&/m�~\p��5)��X����4�	���/�>5KŃX�Iq�̽�0�4��u|���?��ŵ��ԏ�zn������r����Ņ��'�am�J�����*~��E���J�9Q�	J�^Q��J����!0N����>�ڀ���I�:�5���Fn����8��;���_�s{%���TCGz���XB{+42f=�D�*a�R-�X����5��Lu%5�f�'��%�;��BP���'\4*��
{�ʶ���/#\�y�=�i�R���!�)�:��k�\�񐲄#Z���-;c인QNv �R`X\��u"k�j����й�2 �_��PWl�;�ؽ�[�'I?��"^\��d'A�
̰�,��'+�Nz&3(\\�jho�9�6�N���7~�f�)��T�bu\�����µ��YӀC�h�d��
����J��_�}�L��NL�:�@? �(NW#K)��A���c���ὐ��&�M�D�nʁ|w^c��8��˲a�߄��盆��;,6]��S;V�I}�96dâ�������\���DQ(͑���Ժz?z�F��y�1���q�ϼҬrIH3(�E&6���������B�m	E�}3����1�V�;}DMn!��Q��Zs��*��;��GM���� �+1ܗ�}m;%q���f�����&�mG{sS�$��;(Px�"��`?R6/Ey�+�Y�o���
�-yCeeTx��K,�Z��ۖ:ay����y-h��x���ׂ�_䠻�||0K �B��`���J��,�h%�������� .*ٗd�����HSCޕ2�J��`Q�R*E4"|_�q2ܚcI��u�����Ͼy�R=mm�t弄R�k��p�&\��H�L���j�	��X�j}Rtr^��A҄>0r=�N��H�ʢ.����߅Zu �O&l��\*�Z�*��p�u�2	܉�O�IG'�hey�S��C�d��@[�Ĵ���@�����x�&^ *��p�`P}L�Lpݜ�1a��:���^���5��4�U�7 �ٱ����V��d��&f/��<�T>3.��]-0��X��q���B��<����$v́��)�]�!����/:$�p�� �X�)hlq{��c�1[W�J���B&X�S��f�ip\W(w,ꉴ���ݵ3}'�a2�����9u�<c�ٓ��k�����N#��a;�����/��G�Flj7�H@�����Oʘ��ݿ�$����X*ʢX����^b{^镐��#>Ҥ���ٵ&y��?
y�����z�/o'��ԶtU���7��?��I=z���Tw��Br0�W��8�:z�nYWꇉ��_��8�߶���vq�D�&�� AP�#!ZKD���^�{���׾Ų@�о�����l{#�P��\i��>���'p�W(:� 9��(D�� ��sbm*v�<C!�J�a�2]a�=��% kB�So�YWƦ��^[J����w�F�[Iɕ�P7D��Z�+���?�DTŶ�c�B&N9-�$y�%j��lPh�rO�>����4�:W�Ic�"M�M�����gZ�t�8�m�'Uq����$�2\��ИS�'�%��>��&I�#����02Y��������p58������`�n���3Z��Ve���[w�S�?@��d�Y�����=��W?N<m����E����I3�-�Uq�)��*���G|���\H�	i���Q���f�D��WTY�.̱�P��m�ڝ$ه�k.�����_��X8]Se��Ȥ�EÃ�����y�VE�~�=�����/  ��;��c�H�`x�Qŀ�z�3�c\�͚���J��J����Dj���htN����r
�5�P�E�ڒ��?v�o�@�āʵ��\0#�=Ng^�^�"<���+�%r���*!,3*CroN"��"�ɻ��4���e���6j%\c�rM��}�W\E�!$im������BrQǭt
���;g�dY]ڿ2C�D�\�����0��u^�u�Qݵ&�b�������Wd����X��o-F�4�l�+T؝�﬌�k����Lܕ�"f]=N��qATB/0(��G�@��lƄX�[��l��|���{ÐvQ����y�ܧ��,�h"���)�:Jy���,MA��1A�[�����JU�z�EJ�^��[��xG����Z�r�W�}y��Ȁa��i�ﻠ����܍ʙ�I��G�1�w����*�*|AT:3 :�a�!9H���b�f��f�6n��KeA�VT�Ʈ���J �˵�F��H�5��*SY�c�l@����*�<=8P�o�10���G/�"Ax�O`_/Q�NMs�|c��}%���DE��N�Y�����(6�=Z��*F�ȿ��b��߸�S�c*�|�>Z3p�~�˱.�~�>��pE�(	�/E<�p��.9b'dϓO���:���Ra��� I�Q��62���Msaj���Qr�����p���(�҃��:��꒘���ĻY�5V<���^f�~�Q�)��S�^�ҟ���O�i��zQi�(�`������ěCϴ�@r��@�*u��<9곋�n�a�{�1��!���<D����ly՗���b��.�*�c�^��5�]��0��v!fŮ_�+�����?�9��z���B]I�cYMR�\t�	�Q*pB&�<�H�Β��rM,����O�趭?"��$�_�nO�����} ������\�t��䄃=C͞C�q���7�	��Ba`X:d,t�GI�0��͘�Z?Z�9w���H�"��?[�1�(�q����s�#p�Rg���|�T%H�Fb(e>`����9�Q{e��j�=�B��ކO�޹Ri{�j��I��&'-�p)�����c��K����<,��^�ڇ��n���J�yT��+rL[}��/��Yr�U9]*.�V`���8��U�dE�#U���dD@�;�@�o�X���E���9�X�QM��!���	�|wJ$E��(���&�G�s���B�}��� Hr9��sNp�e)��1�o�ӆ��$ ��H�H����>ԍ���#��VˤZ��4Bt�|W�
d�(8X}���#��%���j�8OP�4�����g��j����%0�\�ܡU&vi�8EOJx���R/؄�*�@���[�-�<��,_� 2�=���	�t9���_�Uƅ��ܫ ��.���'�w_/�
QS���|4�d/S������l)1�ꈩ�j���C��[�V��C�|��v�q�Z�r}�/�����&�,��UR�B��5�r�s{�W)	���7.Y��A��:�a�9욅��^��`k��9��B�%����a+�P}:Xr���>Pe�M4 G��f6Zu&�;a.ccU��44�0����eS��Jh5u
�]2{65B�1f�
7d�֒�v�ޜݷtK���a�_��&�%��ȇ�AZ�����Z1��u�ҭ��!+59�2`��Ov@�e5��8�prGn�`c�9�G��e�j�)�2i�(7t*�ϤM����+P\}�Rƞ)4�1~���ˑ�)�Q����V40�L�6������~� Ik ��8�#��$P�G�"Ѹ�y :b�\��M;���8�]5����uSѲ9�gē*#���n���ku˹�&v'��EkK`w�"u�1��7���@�{!h�[������3�eUȥu��9c�b��O�ͫ R�q�E��ֽ���|�`&>g :����-ʩ�|��M5!\��\-zW�7����g��ׇ���#%�#$��Й��G�����`��,����2u/�_J�,�4B��ق�@��g��y�)$0��]����YT����6�ACd� ���'b����)�V���/�/�䊱��of��{"���o"�]'�$��nU_��:�T��|�I?1l��I��y:�Wp@����e\�}�M4AL�3 K  Z��r�"A�d��(�GUWG1X�n��V��0��>y��	
G���)[[ٽF���@Qt��.i-
/�� sj~���I��Za�#�K�-�&�4��{`�^'4(ē_~� ���|���=yS�����2�+�k�/��[N��FOŖ*H�1{|�X��
u�ݕmt@�5�����������]�����\�/ZΪz�r:p�K�$�x�T#!�ۃ�q3Ƀ�����Z�o�=j,Wkl8JS�3��@�k	�ن.�G80Z�J�뎸�n����P�R�s~�A�r�g�,��5�ڇ����)�~dT���u�hx͒$j_m�0����h'�Ö�tzYʐe�u^1^i���Vi��e��ѹA�S�+�ؓ���"��y�~NJ��5N9}`�ˤ�c�=�a.p!�ǳ��Y�����(�Ҝ�ߴ�__�r0`���kQ�����2�ټ�aU9p����+͙���A}����`�����)��D��|�D����e���Q[ģ�q�SgR�4�x�#aˀ�J�ݽ�����SNo1�%��@!U��˛��`�!�aE�k�QL5�@���E�͘��*�gAx��N��+5*�������L���8y4}��7���bc{_�-.���D{7�}d�O�6ؗ��汽d>�:�u�fv�bᡚ��0������w̺�a-���%P��Qn���^������M�’s�ة<���5��s���[7ٽ6��{��:��I����R���I��"��98�d�$���8��8�`:	2A�=Q��=��O1�F�,]�����L�}	+����+b��긦غ���"��=՚��]������BK����M�^�/ЖӿH	�'e`��\�'��}�7�+�d�$_�mijE|Λ6�T�a�� I��ѽ(��
n��e�p����g/�&���cJuqaj��i�C�u�/�E��r�N
�>��c�wS ��}�N������>��j�l?�1C�E�.�wē��F���c�>��k�H�!��;�2:��[�����z
]3��R�E.�ă�f�=�ǻ:�����Zl6*�,���R��^0�����d�Y�䵺#)�f�Q^�:
��=	K��.�}}�>�g�3�G|w�9�}�I�n9�a��M�6�����F��Q;	��9k�!j��Qb}a��t�&���n�D�z�J�1�'�@zZ�mR@��Yr|��ٖ7&'��6Ѕ�N��m���j��*P� #�'�X�g�k���֑�j却
y��Qo%(x"��B@��Vwl]"Vo�%񌋣��qBb�v70d��e�ǣh��,�����+<̖?�^p7ɟ�X)��	{,b�=�����`I���g��.���S+.�c��vs!b�|l�)���P	_~xVw��٘tك�IJ�)BPg �Z"�B�i�˜��b����ՋT4��s��|�N2�x�[���&�۵�p���R�]_?D=h�>�&�u� �b�<�M��j��r���UA��j�gCu��̲�wq��O,&��\4]��d�:�e!��s#"�5��KH5F� �S�f�C�	=W���VI�3ɞ�l�G�DEv��"�����'���=�ŞJah��]�����H�-��Z�t��_*m?�/]�Dg6ݗL-��f{n�' g/v��V���|9HB�$KQ�%c>��?�KoH/^}ڿ�e��^���~/���l ջP،k��ufZ��aW�֚�(D�pO�!hZ���^b���]1(|o��N�e�sR�*W� ݉�ᯫ�*d�A�3܉(e�3���C�{̉ ��$õ�YzIJ��;�3烈]Bi�-�8�~��	I�l+�[���Cl,^�Mܡ��@�����%���y��,�L�a�#�������J)�i,}Z|ղ��`v�iE?;o�`QG��FH�[M�q٠��i���Lz.!��(�@�T.:�39D��ذڈ��b ���uR�Ż�����?�`#밞!����5�v;��%�5S/ HO�L0<1�o@�F'�ô���0Ut
/�>u��b�@V p�`aX��6{�͑�LL�=G��+
rt{rF������c�Eb�����`��x��8�v��E�DB5��1eQ�RO6���� b(�2��h�.MqC���z{�~�o�FV�j0���ny�9��S�E?��F-R��e�������@\QH,)Y��{�4j6�3�-�|�Y
J%�!֣�|?'^}���P��fZ����M����p�XGUH�~ �
���R1����Y[�,��Zڜ�p�*
0��h�'\H���`�3���Ԭnf�x�ŧf������c$��z��ft�T�p���y�E�h�V4�i߫�e��t!��ƨ&&
�&��@0����0(���$Q�ؘ�B���}�/��_�%��!;�1����B�Ăɇ�Ag�N�� ���g8��Y�\�@��
5�x���J��)JT�>�"iJ���8�ךza�J�Uds��Ǐ��lP�3�H��;,r�p����o��Z������-/UY~��|�4[r+W�4V9o��m�ې��A��5�u�v��¤���t������a����)�	ɔ`�m��?̔g��k��_��f%��Ӯ�Q8tW~2�R%���N��a.,>��U�pn��FQ����l�=*U�I��:�֏~��D��Q;}�H�w�[���Z�. ���qTO�]E�,�!������V���i�	c?.]v�*}�m��QG��{Q�f:!(9L�+8�3D���ʐ>�C2t��\(�� Z�SX|z3D�j�^��٦�Ǵ�O-6T�u�X��f'��[x��nV��&%y��	��9%_��p�̗غ�r#y�0|b[��l���Ln������b�qI��0)s ��B�ցʐ ���)�d�4!cD�d)Y��`=��v�w�SZ�T���d%�36=J7�k1-�����ɚHF�LT'B�E��?�՗�df8i	�N���V����Lh�d$�{�����O�f�5Qy���
:F|fG��;�]�m�^�����X]�����E��L�hQ;�Y�����k��a>�X�,�Exy�N���^~m�WU�>Kݡ3���6�$1N��TL0%���t�T��	�,��.V�D����UMs2���x�3>�}���|�{r���:��6��hd�e	����9W��៝�V�?rbB�Ν�`Ȳ\�C�w�}w6z �Ҵ3��r�u�F2�1�yrcA�p�j�g����6���궈ɉ��k��K �԰��)V%�ꄦ��V�.:�q'�21� ��5�uaNT�bwQ�E0���EؠD�q�q;۝��'^��ٚ�`jQܭ��O�t��)�$R5|r=�<�Q��`e,�3��Q�֓p����-�x��7��Q1��âs��p(˿?�&w	6��y�Q��xNS����gwï
���4�6�I�N�
&�@�����:�K�{�{U��cSM��Y��5ނ��eh���Sԭ1��gV�/3b&d�.�&�,c�����Z����Fs��?A�|;�,T�ץ#�&z�`�K�#����.�"�:�gKPn�;�]����b<^�S����z�AC��Ľr1�٦x���Kg�8�K�T4�0>���gj�I�z��'�0Ȃ���K�
$�A��K��MK��ң�_z�ݱ����UN�s���ߗ��AX�Į�p{Ⱥ�����f�"$�$����8�Z��wa���.ᘚ�9�Oo'?z�D����$S�R�Qq�}�;��trÜ!��/���1��^W�6�ԣ�( �cA�)/��� >�Oy��$ưj�r�����5LJ�G����\6Cz��Ȝ��f
9گ��y�u�ϲ�܃P�������3�P�4���8����b�|�bly|0�[5|�<-09����5bbdξ�N4}
���5��C�r��a���mĔ@����t�����UR��+����9}����!�}���T��U�B�(&�-|�ܬ7d�-y�Ʉ��5f%#{�B�D��~ ޥ3��������^j�� ��4�	� �>yA��?7��5����3E3P���r�t��D��g���) �v��Q`B�N�"ǀG{:P�
1*�Vɒ\�9NҁF�paI�)h�e��R*-�h��-4k�!��'׹�T.�֧�A�5LPHrYH�P�Df��2��$����W�co�\)�sm�ђ�Syzx�O�&����I��.H��i�h�!?�&o��p��t����;�>a:�e:�EzWڛzAU�W�N՗�}혖��r��y��t�@��K�RsGy%t�rn؎�`B�.vy��:埛�0mUT���u}��5��_*��W��.!�i���3	��.��(F��CcU}	��Hx^�e�-�M�U9"Om9�U�j����ڶ&@캰e��DS4ٚ�����uo	�rX��{�,s���zP�<x[T��K۞�b�Bc`d��p%:���t��Hq7#m�Z���ee�A�Q͛j�/֛D���A�Ih%�(U��yD���&šAw��Qp���f�)�QUX�٬�ʈ�?Ȋ,}�&�>tP՘%gD�6nm��O9�VZ/5�&�Ƌ:p¼�Q<\�!l[�@I%ufE�~h�|��M��9����M�Sz�ɩ[iY�C�9�<Y>����AB�����hn�R��	ӵ�K��2XC5�`�eGo��X�i��*d� ��1��a��-7��h�=���i(~�c��'ݩ�v�MT5��("K���^՜���',K��O+���Jwյ�����q��_+6�����ي�c�|�}R��&O��/eu�#L����{7)��.���:�� +W GTվ�i�����R������D���j#�5]Ec���ܐ_ށ���_\YX���(�>���Aq�t�!��2�^������&�A���>��KSkq]��[,5t�8�,��R�j��j���!���K@ɢ�`�X�Z���ں�.�>���Z�fѐ��'�*���6~e�?�u{˒j�m��-u/(0��ٍ3����vER�V����%�u��qʾ�r�NJH���c?;�b��%<I�9N�J� .���UZ`n����p�#jS�|�&��KA$�0	�sѽ�:ײQ@ ���=�$���G���b�1QW}�d�)�7���+����0��=�(~2Ku���p��Ţ
H�'\@��xn�k�Y�����l= %bA���>! � �J���R�&?�-�k8܇��E��PS�c�^��*Æ�z�w���3(d|c%��S��#���U(�E�ΘLZvk"�3Q��+իJed���\*��`ڬ��=�zٟ/����]�k�ن�]y�3sV�} �:�#xx�>�.xo+�*`D֟��*�&�J���b��]�6.!�X�c����Ƹg��b�(���J�r�4\9�5�{y��
p�"���jk���;;7�$%�]��?��NL���>���r~�w��أ�afi r(c�X�-/[ĭ���i�rڢe��+c=������xԩ)��I�$��~d�$��OЋ�����NL�/Bg�:E�'�M�03X��1y���Pq�go1���u��W̨�Þlc�4G�Kc ��$)ubb��A4-���dE^����&Ӛa��6�4�H�e��r�d���R7�Y��ol�K�ƻ�$}�����뉽Z�����յ�S�+�Ւ�b|vζ�nڄqʕ����:��g=��8 Փ Ίnbg@�3ߺͻ�w�n=��U"pvp�!�W�D��IK�@�2�D<�`vr�U�e�:��\~]5���T/Z4=�@t��}R�<�q�����7���M{t(��@�Dz��\�$�!�FV��v�vƦ��\XOw���8��)�C��^`��:�?�	Q����o�϶��hU��cq���q{]�?����]bs�q�K�(BT?�>ŗ��������p1�7i�k�W��Nsg�D���vY.r����mH���2C�E�8�7%J��0Ѽ�M�V@gkʶ�}K�\�4�}fs~O4;&KO��nYc���q$����]� D���~�U�,��e�����cƳX�|��U#c�]��8�nw�����p<�/oK�%�C�كͳe`���TA�ө�.�J<��� ��a�F��3Ivx�ۅ�ײL��Ƕ�Mۿ4$�'��8��h 5{�y7����H�
i�5,�UzP.N���F�ݞ�/E+l�L\	1D�>B'� ��_`��~��rCq��,�����6a�K�}I.�4���C}�Zu��'�j g��ׯ�'����37�#NuF�V-L�jtme�z釋#���T�E���O���e7�l�����6�Mq^c����D)��ƅv�ꮱ"���!�I����r�ۤ�z�THf#"����'`唣	���%�Ib@��JX9��;z+����v�!�*�N�p(IfeQ�s�M�u�d�����0��ͣ_�������י��7,5^�=��3��J
;�$l�ш����8=���=��O6+��5���O��Δ�P�><�D�yY�����I`��5rEJ��.�{_�Zh�5��v	<XC'�0��6��6��Ӝ��3���?ӖDd���ř,�� x�O90�P}
��y��.6}�I�$9�c����@ -��R��T��JpL*�g84������ᒅq�#�JkSԼ~�c�%�+��

M�9Z�9��PPih�d�0d x�Y�VLʴ��OpXs�~�5���(� ���fx�M���x+�i��q+��f�ĩ��VH[G��`6֕T#[�rJ�hY%�\�-���Or���D]���4'wQ0��(-�8`G�\�xV�
�x��lh��-eqk�#)�D�I�:#w�o�ԌH�[�)��b��� �K��N��c(8�g�@�㕡�Q�c�*��%(�_��_ï��
�i�d �[�B�n���ڒ ��>e�Q.���S���׏?z�<��䵋�{?�H���c�Ѻ=����7
�8�	��H �nI�!�[Y�����qW�V�HJÜq�����p-:��?�bG�p��1�-	����J�cp�����n߳������]�e����Rq���9aF3x��u���<mN��A.���4����b����;6)��LL��[O3�����<aH���]p��^��4�����02Ac}w�<���~948��, �;���:T?k�apϿ��������|��b�(�-�/���sk>�4�<ϋ!N�p�EM�Q��_�"gԀHp�G�l�������X/�]��PȔ�D_-.�Qi�B��ߘ���S�g�� ��QE�F���а����da�5��W�%��X�U�oi�I���>�-Y͝��A����%��1i!@:Z�}�+��
��c��|A�~oc�����X�F��0'���Y���t�0~ފ%��k